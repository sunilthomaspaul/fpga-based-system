XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��~Z50��##���'���ն�N恨�L7��Q�[c.2%����i�H*�T�M=�M�v�����W�@�&�.7�3�t���c����䰡P[4S S�`R��'"�6�Qy�g%���d�z��%��l����T��rL	6 �LP,5	����<�R��b3<4���J��G�'���r9�j���X�zE���/1=��2�!�}%�9%�1?�՛�uw���Z(A�2m��$I��I���>�Wub���a	C�h�@�%M33��CT.n?~zλ�#�zH�W+��Nl����<�p��|� yI�R�����'�1|���U@c��6���3`g�2l��Ia�p����F�����ګ���Y����܀��ák����SWMx�w�����p!l��0�-b�܍�CE�B!7ʸG���l�w�˗Ů�F���[� 6��f��x��r1�I¾�y�$��S8%�Q�1e��[����'�����̢?�Uh�f��+g�<�ޛ�Le�Y�:��}���E�������\%��vz�tT�\���^�/8ω*w�m�����v�u����hيv��`��O�T��*Ă$o�������A�oc��Py�W;��cC>[kg�Q���h��v�2{ٔ��,�
���MVg;E��1�{9�{�\(�ʚ솺^NG���`�8{�Q(�a�	c�]��5L1���^zt�O?���(����A�z�z��MX�4XlxVHYEB    4564    1270����dw�P��HW�n	�ZE[.\Rpj��Tkhwe]���0\����&1W{/Ų��'9�ث%}y.M�l��2�DZ�ղ�ʹ�&�QJ�������_�	�
����y�K˛ڞ+�i�{�I���{">KCL�	Ф�D~�����A=P'ht3�ejL4B]ϒ+��p���Ri"�X�^�}�l^6��$>�h����!��>.n�E�5y�ULg��������:����tB��z�N�i�b�l�xB�J���f$gg@�׈Bh�}�q��)xh@X�V��	�k��FmTb�u��5l�����:�l�"�MOo�N�J������~݁�y1�$F_���sz�z�id�
�8�`d�� j�**��`Dw���9
R^���<Ș��B��r��\pX�U���G�W�`#��kc�bfe��q<���I��"[�cV�IW� oSp��}�@��&��U��,�@�]$2y�mW�{,�!��xD�l��m��d�΂!��Z�$E����X��/�aT�B���������BÒ_I���ԝۘ����d��T���1�C��e2>���y9!''\�k��NeE�-���
A��,�0�rq�����O��%�:�����F��*�������PQ�噋��n�-`�T ���D������pR8\a:[�;�:P��ɣ.��������+!V�Dl�%0�G}e���ĭm��ɦ��!�=����)�����*B�+c���SN����7,�����߅���"O%���H~ ���� ��+����=F����P�|4�V4p��QM1~eG�r�xg�	h,��S">�A��ƭ�������=Vt1���v{�n��J QΓ��$��"�`=7��"m��<ƨ�C0x�]ɈFZg��|	2W�E��2 2K��]7T]+����p���V�bu�y̪I�{C׍b���r��	�ȩ�#}���hJQ�k�m����5]���3�!.���_4ͨ�9�f�q����\�6V��Ux�))�s�ěM=,߷`^��M�tZ0��^��x� ˾%���U����`�mD��KtFD��A���H�]2�n�B�ܣ���A��/�w��Ig ��訒Y7@�gCb
V�n���� j���C���VI숧.~)��޽��\!�'��tC�ng!�P_Ͼ_���ľ�G�߰1?k�3��)��9xR*x���5�Gα!�o�D�݁������%9��-�,�F���L�SS�_�;,�v��ť2>�L@:�;V��m3���	`��N5k�O�Y3jab��Z��[�[���&$Z"�w<o�֓i��̮�_���u���-T0ĸ���OKw]��rц#>+nuV7d��	7<TS��o��?}�0g�qN��KJ��¦5v��5�8��%�w�ڻ�.zf��|��2O㡟JsMv�BF���*�h�p#N��%�1�ל���w�Fhg�#֡1GW�9�"~{�k��Ǔ$�7��$Bʵ��8�2��:��VS�R�ps��SA����'-�����
��>��Q1�[ }߽]��?ϙ,m��2��-���<`�(��%�C�#����E��*F�4��
��u�f7ߑ:���=���$��j�'f�ƫ_mg�۩��\�������x#�H�}w��[�P�m���9���jP��C�~�?�{�?�Z�^�_{	Oǭ˚�%��)��2�U�����ƙ �jz���O6��-� �L�����TT
r�#��(�<�b{2 yb�PnK9 [K�<����x�]	E�8��ŭ]�I�4�y���t���:��'��Wod�*�G�KP�ag�J� ����^�]���-���1n24fTf���S�2Z���TX���F7��=��I*d�|;7_BE�P��q����߫=׵q|Hh�f��ߋ�]�ffѓN6E�My��_=���`fL-�Z���ٹ�>�j"rz�~�i	�
��_f�Ǒ=��}lš��-��������[�|yd6I5_�ff��'P�����Q�ͬ'i�*�v��`N�2�^�3v�`�A����0���
���^@�MZH�z7$+��ҝ�G�]��\��T+��.�%��KdCj�yXO�.�=�k���|�'�<P}O	$���.x(o�� 	��64����#+6�)x�\5���	S߄��YJ� ��K��z���ez��Yߜa�[�+$�-���:>��hV�E�����Đ��`������Vly��y%DS�䰘ںyȠUJ�	�n���o���k�	b��?�h�%�tb}»����w4ϾΈ�Q�]L6��y`��#Oӟ��i�N_����t�/L��E�L{�.�1��(O���'�)]��#⊕N/9{���l��[Bz������`7����X���o:���U۳������7�H�bI��R�7T~��!���wEא�T�7n��vf�/�[4�J/�'N��lZ�����'�~Ӷ3��~2�X%�8��
�A��M��q�6���.��Vsp~f"~���P�9Y��_)v'��g4ݐ�6��bg�k�� �%shA
GG� w��Vf��{J�c��d���.����e����f��z��Y�ɟ]��Yڒ���cӍ1�`^@�QVi���C�̣�*VB���c���6�c�N�˚UP�җ��|�]�U˅��	5�k��2u#�՞�w猝f�<G��TY �$5A�w����)�-h4�NB0��x�����W����j�V�g=�N�Y����ޜ{L1��BW�K�kO}Xܿ�%����.���-D'~I��ۏ�y.��{�<�ۂ6��0��Uy�,~<R:�3CT�uo��@����&yں�)�3�	 BoBDu�|�'.jP�[j���%���د�G��P _FT����&UjV=�6�bk�!Q�л`��_�Q,LbQ�ûD]#n��}4�Gi��{wJ�uW��6re�c�-e�L�c�7c�_E����*�
\,߄*��\r���m�:�o�_"GG2q+�h�b����s;ɀ;Lυ����i�L`��=��D�̪��Ҁc�Q�j�:(y#�����%4=sZmn�}%q�"��m�L��hƫn�8ҕD{e鈞��?0C�cn���DbA-���H�����>�4-�5At���t��B�������X$f̻�F�U�C]	$�Xw�}?j�g�n��ި���
w�};��e�����~~eH
πIV`��>^�VZS�u��b�}�#t{�٭�\W�dh)��!�[s*���)D�@$c��(�n��/E��şd3!�f�1�,ȉ��t��i�(�D{{�$!�&`�f�U������o}J�84����/U�v!L%Q�~瞮�5��]�"T�����Me3��7��e�y�ť�_X�@��&l	e��CQ�I?�V�|����3U�ۛ�ez����@k�|�cQ֊�v�T�o]��Vyc�uR��W]�Ч�Lc��}��r���
b�sv"0��/�s�����F�����4!	���e(�k�*���A��'��R42�+ѫ�_+����i�o����6U�(���n#(\swVF���%�M\j��]?��z��C	�CUd�`��͠_��\q�b�8���(o�� ��]��"P��V�x�"���?�����'�%'��D{��(�\t?��Y
�Es��_z�b�<fA@dğ�>�>}�o�)��E!������f�U3���(��gvۤeޓO���_\$�`�B<<�q�|U^|�	ۂ�Q�U/ݢ���~����֑҆����^���R��+��m��bN�z���x�T��|�nX�e�se8�
J�8!oM���;��D�TP�>'��|�݉�&>�\���n7�����G�uK-������R��J�*��SZ�Q�����U/0Wܼ�i�蘒�P�xϐ�J�۬�^���y��qb&��	ˡ�)�ސ��ٍ��ݎHS)-�M�rS�y0�365�a�I�.��wB9}��<7"�[�96�d���dt��q�Ы�$�k��+.!L��J���U�6I�g.o���吺��p��Z0���Q]��uq��-�1,�/�RQ>�6��I:Y��g�P���Ls��{i��>7�x;߄��S��x�yd��	�����wY�����f�+��[����h^�GS�̼�'(ncH�wv�:w�X[�I1�a'����<���ɰ#�����d+�#v���d�L,��k�aA����zy���F�e-�|G�p�6�!9��.����}�Xt�l3��m��>,5�ޕ�/�y\.	���܉9J����=u����Z����6��Y�9#Ak�ý�o�?���*��2�9�t�e�TD�j�!d��mYJ�5���� ��]��HJ,C_k������x<��S��_^fM�/m|���y�v��^�މ��I��Zb��[o}`�ĈP��M\��G��l��]��{�#�gã�AMW��O
#i�WZ��n$t�o����ס�N*�����[��<_}W� ?�#,C��Q|�PHk��>VU�su:F�=�+��]�1uDxf�D��.�}��Z���bb85��U1��`�gj�Tz�\