XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��H�m�_(w�\M�`���H��-�˩�~�ȶq���)d���f��k�Jvzx��)[ǜ���U/o��Y�s�R�_D���X{�\�F�ff��\��/|:�"qCո`z:#y)jfHE
� kT�)"�44�#�����oK3�3^�չ,:�w���%��%.7v�q�_�����G��uB��8�`%�;��9GS�#Y����Xɩ��<�¯�4=3��Ie�Żή��*��V�
�F�U��HUso����ވÛ^�wD�~-8@�#X�6�N�VS�x8cd�� 
褶�x�͈Ϋ@�9Ў���~�]D��6�J��R����q�ʷݾ�f�,��ݷ�G��0?P��5l/�9BC���
O��&.[E�Ԉ����z��/kiPF���6Db+lm�
�1tT�EDX�J3w�#Z1n�5�����=� ���L������ܰ�!�YB���֔7A�rAܣ�T�>� �*�(����]+L-�9�BF�G�S�Ns�=��S�K�n�'�q�r�O�&����Y��KͲ׽P��|��j�7牗𼓷�%~��1���ὃ����q��7��\������[����y��p�⛣�S���*K�62Po
��Mȍ¾�9������2x��N���%�q�k��j�.f_�t���Q�S�v�(���]�+\���a0���(ӯ������0_�<�z�%(ʦ��7�M��Qe&��˻	Y�^��2.Un�%E�{�~��yMN��jXlxVHYEB    1d59     8c0��.yx�!��L�Y�+�����G]܄�,�����G�z�OіEِ�c�1���Ы*eb�&-�5��oкzu���ݢ^�s�񦻶<�8#�[�-�����KǊ��|HzBu˺��{���N�j!g����p<�����<02G�8���lV�e<��sh�N�P9��.�S1�i����@W&�1i}��������¼�v�֦r�`#�����~��T�\j�4�r�&��f�Ö��Q	G����f�;�|���o���r�����,8�pĭ�F؛�u/|85��++F!-��nQVa��67)b����HQF��3��_y0	z���P����+�)�E��Oo���h�7Y�Y+�'x�x~z3��B��t9�ѓcu�<���Ϻ�g]�Oq��?$O���Z��"ଜ�Q�����p?��z��0�W7�3x5$�<�G�!$�i��d�y�8a���O���)yUӴCF��G�j5:��l_Ǆ��D�|��z,zg9?�Q��U�Q}Tz��4
p����[�6p\��o�Xʏ�#]���ﬞ��[d���zr��&p���b��kp��<:+��<@������7K��K����:�ɔ�E��u���ࡧY��z%>l��]��3�.��{�Y��Ӽ��ٰ|[�6Ji�n����%�qF��Ą��i]/�7����TJ�;Ml����)=���x���t�|DL.m�KhX±dG-7KՑ� �u?�p�Kܾ���Y�{����2�t9E�pR��@:#�.?�0pG���PM��j��h���.�4�G�Ȥ�Z��,M�� %��W̛ ֆU�ɳ���<�,���'�]#%#������eJe��V
�53�R�G�@�m�z^>*�j���|^�=�	`#�aD��^��-�	����ttip�V���5Ǌ{pn �{���I�1�rɞ���K� 6�u�`V�1��[������_LOI}+O1��ܷ��o����1���ռ�lHMȤOf���*��%�Z�λ�fAi���O����CǷ�Xe���)n�1N�Rt�LTQ��r�>���W��)Ղ���+��d7
u��B�Cf�̓aׄ�P	�7�N���A��H��{��ϫ`h�'�Z���������Z�O�UZ���c
��o��`��Z� ���:�T�ΖU궢�Y_NlA�}��'̧5��u�CW.m�,{B�pYͻ��z�׏��0b����4!�i�Ey>�G�Aq5q8���m��|��{]���X�?Yk]-sL_?S)5��L-ؚW���1�B�:�ݏ��
/��;��0�1�x�qMG��f�U����������<2�j� �����2�
>��H�<ƚ޿N,����:����aI�� ��3�J��ԅ�P��l_��B�n��w�=�7,*����¾Kє�u�ߙcͭ�'��R��,���*ѵ����(�Ņlȗ|u�-�:��\M��bL~�￧�P��oK�OX�����>Y�O��>�x#Bd+H�%S��x��;I���u��
C�늂�$1<�#�W�����MM����
��\-�:���
�����P��A�t �s�(�װ�����q���j7��tr��6IQ�6�
��F�N���l�H�x���c3�\��r�7@�us0JZg�"_02�'y�ӥK�A.0P��nU�>a�e���2� �,W�����r���K��a,�/�u�D�'unp����kϪZvH�a��\O�ł Ík�;fjt�-1Y�"�+�'2Aop��/F6O�e_�Ֆ��k��M�|�DU`x��"� �(���1����)�y����f�����r�*�W=8E��D��qnu�ϫ�����t����V�
��������.s�����rH���q�
c��r��]�]:B��M
U7n\b�A�#	������tL�-L?w�#^u�7QRFF�5T��"�S�x�dtʐeB��t�b����w껂v�|?]_��%���'˱d8XJ�S�{	�*����j�uò2.;�Ϸd�������~�в�%	��^�SS�N[�q��衝�P@T���ƫ[	�E�c<p\���.��iҿ�n�.��gBE1�pΗB��MP��@j��9JҌx����չf�b�D�Xcs��_Qa^�q}�<3A
y�'8}�5A��V��d|:fh1��