XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��4$8Z��g[ѝ��r�H.�
�"�u|B.�S�^�3kx׬B����Ĉnk�J1�Y���Zck"�.z����2�6��V���$R_���8�d����}��*��[?�LZ��������o�SŞ��T�b�չ1:��Z�7|&��!i���5��-6��v�|#
�R<8M}K��l�YQ ���7���F{5�8v3���@7�~�vܸ�K>(S����cezk/ܘY��_��+rF¾�K�[��2���E�F��Z��b�&
�1��&���!P[ԗ\yoh�~�K�/�e]�h�<���������F�VմV�t��oM��h1�֜;M�*���eS�V�]��C��3��ףI��Q)�9�/��݅?�����Gx�C��f�Dm�����h4_`�j
��%��$0L�K��/�N&�m���K�Ӻ���Ok�����Q`ɵ��\�4a�QF��(,�
B{=�������/��N�k�ⴿ�j����$#���g��+g%�ƄW���B>/;�[�sOc�as���_�=��?�x�עb�dFK��f�3H�q�Gil��@��~!"��sA��~��S����}�Ta,='|¸��SZ�Z��(�^d�k^�PVp��1��8��lfa��B����J�vD�b��f�3߿�لѨ2�ExS�x�r=2����3R�9j���'��3(u��/���Hh8J�lc�D!KJ<�O���L����&��3q4��K-��U}U�Ǿ�XlxVHYEB    1a2b     8f0Q|��K|{�m��������F���M��b�$�ٯ[�u� :aZZ�D��SD��kx��� [��-?`ms�����~�����}�]"{þ1�������EZ�o���_�́+;�z	���J����0u*f�"�U�d���I�yb�;AB(�NC�R�K�r�y� v�67&��{h��)8t�u�^-��C	��D���7�A�g��t1������`glQ},���m
��j��h�rE�fK|]Xnf��b�X,��Ba��_K����|q�_��Ӹ_���t�Ͱ@7ǵ(�1������^�3]q2��� 2I��,p�VuFZ�+3�$ҋS��`r��.b����*�P�?�;�.ZK�F�԰�~se����,jVsqk����h ����j��=1��O�n���$��΅�*t��l�םw�}F �:���޾,���R��ǲ����]Y���a���}��#�¢N�1��/�`)�x¬�~�A;�5/ �uD���Ǵ
��������*O��ih��N�X�\Sa�q�{6�Ir��K����(ca���gu��K*Yc?���+(�^��{�v6��ù��WǿTX�j�9��1_� 8�-�i���
&�^�P� P,0[PK��E��[�[�D.�(3�(Z�9�� ����ƅ+�ؚq|���p�-RAvn�}"q�<�u7�1�af7=u�㊔a5強r����_�R_��zjSNM]��*[f�\}�স�O��G��۞]
z/\��i�M��6�]4زI��d�^�<ݔ��[����
8$
2�A8t��w�O��,,�d�w�n�����Pp��E�hG���}�Y�<��.Q�,�P��|��4�M���}Bˑ8��[4a5��%�y��B�}F��m}GЍ}����DY2]k~vը|�J��3�8��H.��ܽ���GF��\�7�!V;�g=�c��mS�����W)w�&�nٲ%U5$�[��Eλ�'�R��+Q��5�5j������?`�(�C�r�ޞ�@��9^��bRJy�����Ov.Ń�1���D�|']j��R�u���0�]{!�x�ӘO|�WឡgF�.vb�u�ߐʫZ��a��)T O���%�`B[�G��p�$��g��j!�	bA ��`�)6ԗ�	_���\�v<b�=]����0g3,mf�<�!�X".� W>�����u�ӓҐ[had�@=�IYz�4���y�d_�F��+���>1���E�Z5�ت�1&����{X/�h*�x\. \O �k����bb�٤�GX����%�n������+8��s)85/4Ǡ�Pk�b`�)�V>/�`x�Q^I��n��FL (gm��B�0�~~K�����>�}O�#�e�l�Q���be�Z� ��ex�/�������e;����1��!Ӹ��ݖiQ!N2D�:�D�f*���Ǵ���$���L��NRw��r�J�J�|>�:*�����Ģ��֛Xd�ʻc	���W6�za7�,`{��_�\��Jp�N�v��鿭a](��+q�Y�E1�LJ21�����gt}/ihi��U�������øٶ�.zY��"<��I͖T�	���?bz�@��`=3�~"�]~8M9��s���	xK�0v繥>=#-��H����H�(m�7Ӟk�U:��_Nlږ��@݋]�ʝ��-���=������b6�"!��bo�0RO���9���S�Y�a��I8�=|Q�z�ϩݿ��~tϰ��r�a��^D����m��~��S��R:�`4|�1��|oh���������.�A�aљ�W�%�=�#�h��/M˳ 
�1��}�zp�#��m_��i�%7u*,G	�irc~�QR����E@K�Z���u�"�C��M��|F�vqB7�ë��C/K��N�4~J'���Xx�ֳ]�e
-e��0zr�����A�yq�Y�<�pA��5�)�+<ۯ�,���j��b7^�,������Uk.:�3��\X�L�l���c��D��s�*���d�[���9�ʖ�끟�e�
/N蝯0�F�t�8���
��K�|3�D���c}"=���*�)�yЕ��R����fGc}��D�8�'|�Chj�t�s%͕��zrc���owÃ4���_�L���9�04�pOcV�.j�uq�#���Ź��*	P҉���
euZ-�\��bk)��i��{I��3�֦F4'%�ϲ�l\��Q.�R
�#
#����2�m�1b����q�,�U����~