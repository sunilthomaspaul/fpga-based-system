XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��#"9F8�p�sv�ܕ�wQ4��3?dq�4eo{��`�K	k}F���2�h��K|nsU!�3T��x�)̝����j+���AU����Ѕ��cm,p�l奙��H�_x��I�v���k�9E�y�������w`nl�>�l�5�F&B��b��{�W�����{��@��4u���8�����J��V�ÿG�}�(򐻪�_�yG�x����[w���٩oGVeҦ�Lfآ�k�=�B&nb���9�N�4v
^�"�E^�����ͫ��g$g�����������v�
0θx ��	�Q���H:���~m&"��T��yN?���T����G��S(�� �?�/�]f���t�q��_���z�%�!��ޏ�6����}bx�����B�/�d�+<�bI���y-��.;��7[QA`���
S��ݐcF,�m�x�^�Nh�սP-��o����+�hyF�����k.�)V���l<A��܅��Z��xYJ�����d��s4f�yZy�޺K��'��+>#�C�Yd��(˚�-Wy�W�"a2t�v��D|��oay�<�B��-c`W�7s��W6�wQ��3��@�Xr�����[ب-��J5� �ns��Xy#�Tؐ玾��V͑ze�1:���Ȳ�Kϻ�f����86�\�L0�lX�nK :�&�ks~@���-9d�L�/?�Bo�p��?bxNDK�t��m�DH�6�U�׬M����Z�5��n�I�IԈ��JWXlxVHYEB    bc57    27e0���nܱ���"��M�����P�S�i��KE���l⃎���@k��@IHy�
��y�(�Bqs�r�!��`�r�s�	[�7lmj7���������=b���{�q����1/$PP�7��KPF[k�����Ϭ��IYaH6Q*pm�b�
+�z62�z�\Ǵ1v��'{��s;�HJl���$�=a�SN�7�RPs.�M
�j�~��7G�����b�5�!Vd�Rfھ�ȿ8
C���tg�Ut=�~Qԋ�T��-.ޠ9M\�2P�k	������OeUT�2�T�I�k��ז2�+ܻ)~r�����mr�~���,L�%E�#>DQ�]f�`�ne=9�w�v᭑j���yI\��;1+6�i���?E�Y\b����x�q����yv� ��̴>6@˘Ӓ_U��=�ũ����Ǯ�P7���Zz��
��KZ���}�����QY2��N�R�M�h��ղ��Ns�QyKu|����#�d�d��ǲ���!@�KY,R�5��[���E�l�� �C"<��(�Mu6�\���⣇K�	��k�Lt���Ҍ�"����+՘'W1=ǐ2�w�ІNZ|�0�yٙ"+�7_t*	�����PlE΋�Ο�ː:N�#�1��K�R���%GG
ȟ����}.O�~(
�H�Pt�&�
 @I|Ի�������b�l@�9�*���Bb�d�K<�Q>����TP��Z�
 p8�	S�o�M��3�C�A;��.V����|^7�Ά��N�V����@����ϤkO.�c	�\#<j�\$��r3Ʀ\�]�:_����+ <�صN*��]ǃ�qT�<������U�t
T.S$����<K|�@�w�]K��]Y��l�TOFx^nԤt/�9�d�W+�8�輔�M�Z�}�tn���{dD��5@��JWD�".'����Br��Np���J,�R�ƞ�Cc>��Q Cˆ:����:�l���#2*՘-Y���6�N�.���:�� ����Ӟ�#�������wi�>�.��!��Aا]t�ᠺ�8"���ag�I���;Eab�l='va�W�͂A �Êb���y,Gҭ�������4��E��.8���/U�gN��Wi��"�K�ʓ=�1C�!��y*�5*��r1�����2TĎJ��m3Ⱥ:-�_���\���v����YugX�+!�B�R(����%�N���^
1b��
3��YQ >��=^( ��Yf���#Я����9k{�!�Z�ci��U|c��"��v�� �h�N���� (��o_Вi�~�6�1����t�)����RSq��bXRrUy��U����$XV6XgW�oc<a��K<���F;9U�q���ō�6��8`P��ڋ���{�B���-�*�&Z|���i�/�Q�?v��{��-��}��O�PWo�$��x�j�<��K�on4�`���IZ��TGq���p2'X�-����x@��ZP��X�{b�\m�X_���Jo��G1ͶS�$�t�3e�URRMԹX��Bkp���E!�"0����h./eh^Q��u�2�1/��C�nHI�œ@�'%y��W��J�<��/|�c`'*tP���[�]@{�I�ʜM$I�|ɏ��8���xQ�0�����9��LF�gm��lZ	�/���� ���L��V�y"�wm�e�eW^Ư0|���i��l_�F���U"��y������"1������&7���݈֩��`sm:Q}a�1�M��Q�F9j������$�F+�-��O|�'��Lm�.�^�I����x�,�=4���t[]�h���?���`��NV]�&�VE���p��«z�ߞ� ��ê#���C7*�g[���N�qJ��������Ѭ|]�͌��KU������dm��=��p�)0� �@s��q�d�k�!ܜ��EK��JS%�.b�E�����Iqܮ�Ӱ���8P��/靚8�jk�u߁�O*}���wLRڭ��|n.��=��'+�oɷ��4��hG|'�F_�y�R�S�?��.�]���E�-��bIo:���M��:��$|��8F�CizhO�PXZ��%����Yd���Y;%t�m:�/T�rJ�a�?�	�Kn�AM��Tݺ��Wz�o��6;��\Z��..)X�w�`��/��{H^����"��6�*c��S���P��I�q�y�"��s�J�Ͱ�t�����lE�;\j
Nw�7����Ӷޏ��ғ(Gܖ���e���I�#9t;��)�' ��%N>�K��_���lm���TM������X�r]�\�%^m�צ+iݝ�I�����6��T�գ!����dW�{?����K�#Jz�kB� ���MɎ��{���rX��>�� m5��
�C]#���/�6qr�����Ǭ+=���x��I���X!�����b���dĩ2��q�e��n��|���oW�n* A�O�o�)�v�1$�Bp��@��!�%�QE��$:���!]6u9E����@�1Dz�T!@Q�+���dHR4:�b6��*������@���<���\�˵bY��l$,c)v=��!��).hPU�������2�Cǲ�/�;�7Pw����z#|sZ/'L�E�3&��1@�`*L�����%��3�,t��PՃ=|���R 0ګ�ڧ#�Ü������[�5
���-Ei�?�4�4�H��������@��lDx:	�5O��y�E���Ǻ�u�J߄K��T����`U"���pHO�V�$��A
�L(��)l��t(�\P���l�&X����u��8+���޽��$�ңK�gz�`�
-��H'v�X�*�s�n��m�30J�G%J��
!�b.�a���=i̻>g�����9�����F���J_��^d&�|&`IɌ:�C�zE^��l)ݪ�l�C��da�}�v�}�5A��Ŭ�ǔH^+�̝���"Cs�p
���g#� �s�ZINj�TZ��Ab��[��lB8����Z��d�-4r��tى��[h5�a����$y�k鞮�آ�TM��	�}y�ȏ�F�;Ծ����{��K�����I��cà_3��c'�3�~��͚HX��v@/�z��K�x0J	4�B)8��˺Uu�����{I��T���9 �Q��Ѿ��v���S����+˂MV����rG�=�'2$���~��A��]�,��`������g8���hWtk���+`�UΛk��U��}��A���~.�@��ٴw�1s�\��4kq�)��
��r�#J��t?rC�2Q��M�ᒅ��
�O�
�8�tA�z�l;0^���tpo:T����/@� VY�4N�}c!Z����+���hĈu錛��o�@�\�na���������)��$�k�)�s�X�ib�yL<�3nj�*�5<�#V_c�q��>ăY�ö����F^�Aȼ�~Vю����.��D���ef�E�J2��@t0o.a�c����Q~1�ʉh�'(}�R��l�m]���
<bd|�I�� ����EQ�����8�-Te��]����6"d�ro6��=.z
l�(x���u��O���_��U��j9]��G��R�tƣ�:7���$�<.���_�Qr[�a��y��T�o��b��ǪH��FH7'��ٍ?��b��kϰ�ӯ����
R �K3�.���]���#s>���&�/W��\	�6U��rhLf��M�QY��{`�r�P��H?�"�Գ}&;� �9E�S��{Z
����=W�O���k�J+�
b|�������ԅ�o�p��d�H:gZ�0�9Xnb��-���2v���k�W���f=5�r�p���W���a�;<�����g�\�E�J��h�P�І�%�"Ub���f���g /����#�=+��Yi`��]���err���O�x#���u3�8���H����� 
R���7��Oc��e�P�e�]n�.���4�{�,�Uԥq׷L�Ԗ�� �%�\x z�7`i�ňp�y{m�0�|]���i�����X�o�j��+X@�on�;b�o���2�*!5f�ܼ]SsC�O�'n���OQ����W�C�p��y-�T�\]���u�-M*nBLzdĽm��|�XڂI�Z%D��S1��/eTH�����2-��X�e��:2\x��ݼ×���������:Ns�y��G�m���ta/�����O�P!�֦Ӷ���)̹J��#�;��0����̓�bw1��kDF.�����C����yӱ��!��V�z��#�q��z"���"�_�O5�H}Y'r8��d1�"�͑Sk[��f���Q�9���}��$�q8�RZ-�$�&�R�k<�C�2��gȬ3?�H�M�)�U��z{�Y�a���ht�ˊ���G0+�}'U��K�ܪCR�?�����|�2�lĳ2��H>��hC���~�;����}T����(C3�@�B���j�p�_h/��O�W� ��wؑ����R���&ى��$o���7[{��iݦOI�7�k�zדx��&��)t��ܬ��_9,��'�q��ҧV�;Bɻ?/'b�*�1D�Aj�sPzG�V�I��f͓�8�o�v�1��q�����.�?�[s�I�7�}��;OM�4�Ƨ�� ���,3�����&L8N���	��@�6�dH�����b��+�=�t�g��GS�R���JxF������1y&��O�����S��"N"�Cp�-���RXc*d Ң�ՕADK�"}tqX�pW�Yr��	J�!��7K�7���q��"�:p�����"�	a>'�����4ml�y��,SDv[I6d��qAvs�r�5���<.Xg*dQ��@�ss�-���}��@R� 1_�|�^G`�\2��]��u��0o�:��ɢ���8,��ѓ���<O)@�wm��9��� #$bc̢�c�f�AEw�zN��jԒ��t�W����5΂`����|���]�iV=&������h�cp������c<A���L-.V
�<\ԂSqڟ�|w~X��\��s��/r�4d,��V0	��h�3"v���/6��le\�MĜ��2���#9y5�����v��H6d�� �) ��D�*����9|��������Ы��M�C��3��Z:un�tz��,��W��צ����8�a��Jn:�;5w�A�����T�(�J�����'۵?�j�Ȧ��U��6ٌ��'����B3�%�/���UӴf1"\Qt	­,�I
��l.���)GN��?�,��E�=��(����Ԏ�3���t��1a���5|��숇$����!��&30��&l���#�i��(��P:�>����" �8����}Kz�nI���ʁ@�ˆO�J2�w�hj�� �J%�t-����~&Q�h��ag���>X���$:T
������5L��&w6�X��;p5%n��Ƕ~uV���`_��bJo`�W�9����THE8r��z�f-4"5�k�h?C ��[+\b��{�$�6:F�x��k�ny�\rj�O.d}2�D�0��������ҡw�OS^�0W����Z�S$�FUp�Q-�"��0|���~5��e�x)7��Q^��dHB�-�U��(O{>ĮC�%)3�,���o���cH"r���gߟ�����;�u������a8��/gbj�>��
�˃pk��U���s߃}&b���ǅ�4��k"'���-\�O僘zpc��9�h����p���_X�>����5!u�;v��U�x�@�������bZ���Dn��2 ��q��%G#�VÔ�X;�@.��f�V�5�T��(�k1���3P=H{v�Z��Q��r��G����q�K�#)^9�a�������n��UKBП8y1���$�E/�lw��6�0��&	�&DjM9:(�`�. �S�fex�7��$n��ߚ}����3�ӽ`�&��7.�L>�	�۵U�\��[�"�r3}5��K���ħ5�mIw	�c�^��\����y�?Y~<g/���&J&�A�j�e���#���gT>��[=�&�k���K'h�����@Q�y2^"%K��1��������$�ގI�2x&�Lyd�Y�@�k��(��ʟ#(5+����b5mo&��.M�'y�7�	��e�����>��.ʎ��Q����H���N���3/18�f'��� 3��f�&Ԁ��=-Í�G��+���l�!|J>Kƨ?1�-e��d�U $(cx[H��/�lm�ʙ�5�㭿W+��Z����t�ءE!n��p�˵������`H�Vl���0g3�M�phW���hT���m��9�����0H����^_��Qؤx+X��*F�1���ڄnͬQ��L	75toC�N��<E��ĳ���g����$�tUG�;8�ڶ�=30�@���d ��U��d.�e)ڛ�69�-N��{��q拊�,\�|�9��ג����>hI�լ�(�#,ܩ���o�Q���'P�TɏZ��涥�{�I��Z?�����;SW5��#��l�E�nDk0�Q��P� XN��斌�_��%�24>j�7`���&<|�ߞ&��Q^Y᥊,R1�ӑ��.�{Ol�%���W������5Ss���x��{���>�,�C�<,P���0�+V�W���� X��ӝP�wBR8D�ϩ��/��R�� �,8(�G�>x�}��Z^	�3��3v��A��3U����g`�vfF27�7òk�j�������&�7���9Ka'��� Z�jQn.���h�� �O����r�7L8Gy���˳X:����C^�#<hz^�S���Qs�m��zȚV.
�e������&�y��>� �Xu�צ���=�%��K�a)f?��\:μ���k����!1a�Lb��W�Uk�����{��E����4�{��Â�џ&ԙ�^���~r۞��h��~���@����>�������*�9��nm-.˻�s���N��'�y�W����5� ���7�E���ٖ����V��<�ŋ�0��Ƌ��#�7����l���T�����!9��������z�Q@p臮�!r4�azu�����?6����n�������l�8�����T�Ѓ,�
�C�,�������	�;o�F�W+�,;�vf9D�ţK﯇�����6�����1�h��`�(���M�*y������<�Ɵ_��-͖C$���{�$P�=���%f c	��J���J6爒ʰiԣA	�`2�%�P J���	V0���x\ěB�z�_��^-�2��1� �=�^�r<+�Q+J�����/U~����%����+���D~k�k�Ԅvv��o�Gy�rw	���ZڥQ���-��b��F0��R��`q^6�V�[�n�N"ȇ�ҭ���]�Z���D���C���;�`�62�O���+�R�i�c�y'�%dbĭ:�M���"~�����N�@-�p�l����S��P��HDEu��f`c/s�r��bꂚ)��9]4�"��5�~�3Gi1�9L�Q�)��I����ȇ�{
���?���O��EdQ�щ���p~�:ea�R>E5�C���mu
lS�k�f�Ym��O<����ـ1KE^-�Zl:�$��hb>��@	,Y"?}v�4g>����7_���vo-rNH,Q����[��	Y�`�W�M�<�� !#T܂򣍘��r�V��<�M���띅9QrKy��_�E�����ap8�4;	��c�y��v���8)���'H� 
i�)۬싉��k�/� �o9�����F���<�U*la�S�`�!
/4���>,�z�PVa6`�㳾XF����N@�C?�{C�>����q�a��xЛ��I��S�Y��(5�d^�e�����P�m�Qq%-�?}�2��q|��C��ޮ�1��)r^0�G �n;զm�%�+kƩ"�]��ZE8��Νh(&i�Ϙ��Cnx�~�����)Q/|�6e��^�@�)S�B��d�	���W��([�1�?�POs�u~*(�H�Ӕ��h8�$�d}e似/��R� ����}Gp��Ӥ<+�\�^���+�Fk�SW�ﮨ�A"�׈Z^��:�y���^�l,^���W���	��-*���a'���}�;����ſ��m�X]����e��e����8���z��1X�-�Õ ���ݷ��������7��|�4r���ȑ���L��,�O���T��pC�����\�Sϡ������d��S��wӣ�oeLK;���`#Cv���x`KWj��E1�
�c��ڃ��=(k�ΪP|^�꒶��d# ����$�'��)d���ىc'��ςg`�HP�NZ;��6�%A�L�gN����)�I�E�a���Ѹ��qf�I ��]�2�����&W���!��߂:Q��g�W��ǵ�C ��Y�����~�,op|�B�%�S�l��SҜ��jb��=>$%��P�O|�)�TA�С���`ӝV�XR���]�dLkm�@GN��)I����������4g>�9����4`�L���O�����Q��X�h��Por�&c����¡eg�$h'�����%P������u��$��Da
f���N�]�)��M���>��)�A<qBW�V��V6��z��lK�@b��ԅ��y�"��Dպ�B}�c|+�ђ����8��e:t���>����$Aκ�D�8j&[�-1ε��5��c|���$[�ݡ����k�S��UΕ�6'#�ŠNď��(75�d{��;��Q�����@"â���l��T��ܖ@'���ք3�_��s8�q�w�p�*�i��o��r���0g�J�x=��Z*c2�r�r���V!�$?�E<��8�f��,�o��E���	 p]�5�K�$2�w�:"�Ϛ�q��}��
I\�D�Q
���S7�_� Y�+�0����Y�Io��r	��e�-�l�|7�^R0��:���nM';[�����?`���o������ͼ�2xm+�eYP���_���!G��k��@����
���������y�pua�N�\���r��ч����)�U��Ĳۻ޴)�N|�S2�J���Zz�3.�{��2�ݍIƏO�E��%1����F�B�� e���~����تF��&��+)	� �>�uU��X�?��]q�O֙��5��L�͕|qp0iۮh��	F�R�+��	��A���LLpp�\�zl����������b{�a$�=��%{�!�������G����A�䴤,�+|��Y2�CA��6�T���U�n�`���ǒ�)>�J��o1��"}z�_��NY�� ��z�30��q!���4ީ*f&	c]0������Y6ȃ���,3<�egT�}�pxax��0��O,Dv��C����bC�b^������)x{_�iߊ\�)�a�7E��g��pl4��=�H?Z�ao�C��`��x���D�����o6��0�vS�N#�H��?5�)�s6�6<�~ͩՄt��o}�8M
��m�;�.BE�&�H-q�uWd1Y;�ȵV�a޹&�w��"�v#ď0��`5����HP�� <	�`glk���i�2��- ?���5_Vݕ�V�j��T��KG颕��?�x�m���*�����o
s�� ��r��AV�8�:���w+��8� �|�.���<рw�b��:��ލ�v�rN�69g�¤	Z;Ŝ�G8 �o{��(�]�+�*��~�Y'����m��|����G �@�g0ݹ��].2�#'~�fx�M_I�ح;44�=��h��{���O��Ei�@��s��]n�u��)9:��Yrc_�r5g�ef+pGd����:X�0�m5��ӏ\1/��k��ҫ�ylG��X:�"����P���x�m��ӄT�j_�%g�����cф�X���ﴇ�+Y���Қ.��`Gz���a6#IvJ�z���JNs��D�Ȼ�y�K<