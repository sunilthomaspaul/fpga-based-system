XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����=��)�	��L�n�����
���xxB_�/�9f�b~���I��Z6��j�� m�f� ��+�}~�e�.m-k�����)�,0�4��}��s �`UU���V��k�w��7g��0�s����g�R�����Lޒr"�c�[`��{\k��U�/-�����<ā���ǩ�Z������I��'���Px����`O"Z6l��]�э�t�kX�dx��1�2j���6!�*�B��Z�����NPí|��J�#(9/q#3�U�����6�������f(Ku=X��<�r��t�lsʟ��S:e�Z����	�5���63W^��4�р��q��r���G������ܩH�鳞)�צ62�5�r�QɪQ! ?�	�m��ᎃ@�Kf:�<Ђ���]�(���VSz�@p8�R�"`Q�6��n?耸�ņQ�=����簞��y�H�Z�yD�.�Qhj�3�>Չ!��I?��)Ql�ݧ�]zJ�+�|�r�l�Ή��6zEe�2�S|�{�ދ2��a�����{_m�O6զ��7�0�hY���f4X�����y�hyo�u���=x�4S��x#��s؊���G9��e��Z��- u���aӈ*;-��]���$՛�Ix��6��F��:C���7���H-z�oR�7\�����D�/Ql�$��r�஧�����+L�R��~5�m��}����}�v�IH�Xa��j;��R���D�1��#��2�d��gd�F��Y$r�a��XlxVHYEB    1d01     a20]����9��	���2-*��`�+��j�B4�1����C�M �zݯ���#tA�[�
��'���7�����j�k���̌��^Я�a8\ᱜ�Q��p��1	�R���ʏ���7���Q1q����l7�7#H��p/��=h�-�`t�����v��˙�<�ܗe�)C����(���e��J��R�r���a��Ʌ��$�&�����&�7)^���Ej�,,X�D���B&�/>}�f�" ��6�O9ɚd�+LŴk�ծ�`��U
G��y�Su�o>BW��%	CGj
��7�ǕP8e��D�o�S�i�"m��&�N�2�������av=M�r�%7=KV�y��j�g�Y��B��W�5eC�m�=���g�8e>=�����b�GZ�^�ҵ7�U�u%Σ�r� �!VG��V�!�Y�bT臶."�5�l˃a&��������Og�N���!� H���C�)3
8x����3z.��&������w�aw�iC28���l�+�Mw��EO��g3�5]Dȭ��(��g�p��O��݅� �����r��1J6Fo)2����N������qvKZ{/X��\�fm�T]mʶ��9�����!�<���R�ј;�uQ��eO�*"���� W<H'�s����º�]f�H�e�����ҏ1�n�-�r��5Q���0����w'L7�į�N���P:?�\�K@"ʎ �
8n��˹/]����ٿ�FX�sI}&h��E��W���S8J���I�����εQ��%���/����M���X�KW�-xz4�<�ga�Z�{��_p����q]��X��]����jTZ+ú�d("`�.�'���f�GK��6��6��.��x�\9�Ӏ�t��۶Q���~}/ȷ�,n⥄�K0\�T�qFN�+��O���$��P�<��+hqJb�t���i �)vƢ�J�g5��/>7����llM%F�Q˂J@s�1w�xH�5� �z'�� ��א�L�99'<(Z�.C��4}��d��1&r1�����Ռ�u���)��D�?�4���r̚]S��D��q!��s݅31���M�	hÇ�������r%B�1W����`�]�B�g&���0a��7��j�&J����z2�89��EB��G��ځ����3�i�QX4�6+sg�&mn���'F	���௫b��o���6D�lf�������b��!.~�����\a �������|� ���n'��=,�p%nPB^�+�!5����Y�	D�(�-��W�\���B#�>h(a�%"ll�KZ�T�X�qǗW��O}�z��*�6���{3UE�&p�i�@o���տ���O��H�W!��8�=k/^��b��g��O ��BJof���J���HL��ȍ词������ץRG�A���ƟWj��pI��3�R�f��k}o���"MK\f�)��}�r �wZ���
P;���]�yD��3IE|�\+.��eI(�!!q���!�E�n��	�fB�oZ�FQ��̌~��9�M^(7��bs&�v�G�3#0���F����7qF��C�$_��������	�!����s��̴���a+�n��Ԩ(��3�
��NF�>��p9��4������*�I��j��VX)BF������g�p�T'��s�O!�6Tc�	2S	�?~j������6��ō:������%���DR�RW�:\�g�x?�E���-�وW�Gy���r`�u
��:��vr�� ���){���{������z��g��Dc]��1��_��HLOb<�B,����S�/�y��� �ac�{�Dp�V�R2=z��*��L�(�D����t�Iْ��e��-,l���\�D-��k����E��i������°�.]�ZV3y���	-��a���l�E����ľ�.���F��..֦3O^����i4^"��O��\OB`������{��g�< ���|�.J�o����<?M ���B��� � �|#�u/^.�op۸�,���m�c$W�j�k�#�d���lj{(�T�Ohu;��q��\p�>���1p\�jۋ���u<���F��()�}Ml�2�r�&��'�����9�t��j>c��Z�p���s{���t���F���,�r���z��d�aDO ɺ9<�'��$p�~�>�=c�oj��z��ߝ�)+Dd���|���:}�� 4�*Q��hc�3ō�݊��`Np�u���G��*9��䀃��|%�b�zY�]�b�J^PoB٘)l�l��Y��u�$�1AM����^y�֣U��s�h�LJ�H",��RV��-p��	�F3��+��~��� �T�4�q�4��ih���eF������u\�D�AԶ�U�Iz$�ݟ���聳^���)2�6!$����F���������TN��]����S_����W75Cɵ�Ƚ���q���u��P9ra��%[��ZN��c+ɒ���^ ��3vaM�l�B9ّ��