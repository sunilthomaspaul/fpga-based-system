XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����8��\��\��§�vD���k��΢A �w ����t�����a�R}(1FI�������&���9��E�vZҫdC�������W���
$z����K5Ld��=�M.�ԁ�HKv\M�?���L0+�֫�QEy�+<q��b���Ch�_�u�}\y�@{@� �Qj�Z��P'D,�����r³�eo�"˅ѫd�.`���1`�7�D$�SU�"��P�~�Z�����O���YR�fϕ�tT���q�n^$_�Hݺi$Jj��`'�Lb��.��5��l��pN�reQ����%�/N��;D�tb�I.�D��1`��4Tk�� "hB(�9-���m	���� $w��T�\h{(y��Au?��@�خ�!w���`1�ر�?����@��V:K��rNOs����ZW��g~�|�a��Ϫ�2�A����ʻOv.�J~6�@�� Q�S�b��E>�������^zht���f��M��=H,clVt���$��3��[&�?s&�	 �#��S��[�y����R����}�qnMEI��[�Q�-\��b�ҕ{~�$�Y���<�U�
*¼�i%c�DF�����=�����}���7�sK^!!��H(���'�f#��j^�dnNM���bt�#w��qCژ�� �gNS��̴x�Lşb�@C���'�O�q�U9�㽑b�o5,֗�hV]��(��7Lǖ��
�$���|G��%��;�u�{<�6f���#,���'�U��-��`a�Q�XlxVHYEB    fa00    2620<0�у~C1��*���#��5�&�8�DNM���ӧ�-���O39��u5U�w}l]S��^�mT�k
�kO��R�Բ������y�x����̳�H��������S{t�����x��C��=�|���B�~S%w�"�h	qL6���Y֖&�N3��K�ˁ�o�i�{��O̮��q0�<��T:�xx���i�#��?��7�,NN9���Yc��5�i%	gJX¢<��	u"�1#38����Sxd~��=B0:����}G���E��<�YA�4���q�����0����}Ѱq^C��C%BVH�xc���gֳ�[��?6e����i�}�XV���K��<�i|H�,�,�F��]~��X'����y��#si�SY�S&s�߽L����P|���.���	�ʡ]bd��2چh��xGF`a�3��F�Q��+���^C�O�y�����l:� dj���'h����7B��_�v���
�~��1r)-���F���!:����ހm�9[ ګ�%�+"�����V����^Q����)���.�h�n�M������5��m�΅�S
�ZU}¬��GC\%��`M@��b@C�mΝ�Wy�8��7ݲ֦�,a ���m��R@?�lh7d�n��\.�e.p�0�{����v"��� �����4o�?"�t��:ĝq���5�!/a��&o����s��9t_�Α�FK!�ah����_|�u�0]2<��J��Y�k�%7���|�v���z���
ȉ�Ѩ�,
V�+�Y7������9�;��"��X��v�N�������r4Vo�'z���F�)z��K�
���RGȂ[��C承Ԃmgt�s=)v�2BÂgƵ�u�W�l�(B9*A�J�~ `����/+j))hT���� J�?TY�x#��(������[Z��)�qm_�^�>Efz��gh�T�7B�S$�WN!�K�:۠��5^�ʯj�ײ���S������x�m��V�PDo\@��h�pdcĠ)U�@d�������G���͚yx��_��cl{M_�?�v����-���·tV���vU��&  �5
�z������=��\���^i][���i��,m߱�w��qh���]ﯔ��ؕ3�g��$�%�%��.6<��_�]|	�M�0�����h6ʾ*��Y�G��
�9�M��j�S�P��-u�[�:�ֲ*��Xڿ�q�_��Yk��t9���Q \�^��2��\w�h.�*��>ANeYX/�fVy)@�N�R�:!�ܔ��X�\��ޔ;��ِw댌C[��σ[$tW�b�t0��#��WM���*al����"��Bd�4j�e��Ï��^H�O�E�9�;��dK!����T���{ 9E\GN�3�A]W)��×�q�F�A�f���QwL�R�>D�����|��d�E+~��wަ��[yY]�#���%�h6��FEi(Q���p3b7�?'Q���zS�wx�_ĥ�L�ꅮZF���_-���s��Ϗ��h(Q���r��~������`�`cP��|��k$�IW�#Hd<�]����e���Gok�J+������eA-�7�m�$��)�ź�}��&^ :�c����r���~�.�T\�����RD��]�C�|:�V�]<��u�Gߘ
EE0/�.(�9X��
���~og:w~�@(�@���7�c��n��~yb�L����4�9�J*)��78O/Nơ��r	����?���U��+u}�7�M�R����z�D�~^��!�n,{��2��-��j\��V�;��)����MB��ux1�DK��לW�d�w����:�|m� �<L�]�+�'��R�z����ҽ��^@{��$�U��q �b�����lf��\i��|�@�~��j��d:�tј���S�r���a5p٢� '�|ᵺO0^3Û�R\��#Y�b�qaM�G��<*RZUd��h��3m�b��͂��;[H�.�'��F|=[ �h&��m��ίօ��0w��.��GS��~��2/H�Yt1�R�?�/����KKc!�B��*�^��C!���ۆ����	K:�|i����LrGݖ���UhN�������_(�0W�`�/���Ć�Z� /�_~y��\�0O ���C'�5�c<��l7���.�a��,>�^K��}R6���Y�Afj�j�Y7|N��T� �Xq����s�!v���ڱj�E�|��!]�	����*z�3.|"���P����P�@�R�)�<�^�+����A�v����.y�s�b�5���xH�l��~3�)�8fk0W��)�g���<2�p�壚�u�y��P����@�3����D�ͮ�Z1�R�%���b�7,5n�(4! �8Q8�L���,�ŉ���g7+� �����8����N��W;jԶ/���u�uZ�Į6 �L�����e����u�z��O5��=2�Fࠗ��
|BI� �G��5A��7=�b!���%��ʺ  �v� .WE��Q�BI1筛e�/½f~0��?��,?�̄����J
S#��w��G�3�Q�e�����y��m�x���Vq�~��N��$k���R[�)���f�?�ӓF���U�<���C�?\�Q~? `2�c�Ὢ�MzSf�Gr�9����"�^ր#�L#�6���%���^6r�F�j�$��;�H�WdS$�.iV���T��S�Y�M�p�0�%���~D�ƃ��]rv ��]K,�`}�5��rCl��|L��U�,�Nw1O*>�;��V��;�E$�p����ҏZ�S�<k�܆����e�����	��?<��u!��9��6�J�TL5=��I�.2�膣a]��1̃Nt����S��̚���=��@���zk���nםD�zX��T�,�(K 
;���D�a��w������>7�U�a�dtL4w�T/!O�-��|F������K�[�L
������ܛ$�O�=�i*$眬�L��k��N>y4���#Lw&�B�%���|k�ѭ!��h�E���]XWC�f����a��`��SU�v3�-�0����s^v���X�6�u�sd�`i��S��*�d����O)��pε��g�%$a��:3�@�p"=��6�{��F2��e=�'?��]}I� w+>�d�t�L��1����/e?�mD+`�`g��~S���D�@۹@AG΄ln��Q��$}����ܪ|��*K;֍T����?�'�	��K�I�+��H	���u�*C��q�Oc�����V
���o�Ċ5$q��v{�%�\�e�휟_��Z���5a�&ux:%Nn���B�`��� ��z,�}��h{,R�MB3���V�0+~�%4�5~�6|%�!�B�|�u�����w4F��B��P U��'��A��/�N_�����F�Ѱĺ�EI��U�������4�Ř~�Y����[z�@�"��*�U%:3���8��AԯG.��\!8��c�F�3���Z?���2
|������q�/�l�F��U�Z�`�G� m�~oO�3ݹl���i�t�*a�k�	tD�!ȢϏ��8�Ӓ�]Z=�E��ƚ�����������ުf������c�G��ni���H1k�K��@JO�G��W�Dp\������7R<�|Ȁr�YE�28�к(�l��U��p���e��Y(�����qġuf��Y|n�����ܖ7���4��{�_m{��dnQD�;�Nh�m�R�sym���w�Ѹ�TM��ͷ� �!����N�9�_�h���d^�������*��SmY����w��� ͤ�M�@��ŷ|�{}[Qs�Fo�#�(�Áb��M�B�+F̕����Т�08{�*T��}һ|0�(��m���/�RP�∯�����L��ݖ��/ؕi��=zξT�pR�j%6A���e�&ν-ޔG���1�H#��\�Ybв���eZ�
��v�`a���.��Zzl����0�P[��^zw����
�+�(k�ZY5k��*I��˧�hP��#���ci
��
��i��Ew�N����zۖ?|���Ub�/�cY�ى��2Ǧ�����/��1��x����Z�m��¹�anwm3̸���F��*v=b�P����]$�G�����f�5� *t�v����Mu��2�|7(�ۦ�42n�y:>�wz"Vv�|�y�7�u4�p?��'$]W�$��(rw�A���������۾:[��+�����v�G����PM=��/�J��^�A��G#�ҎI�8$|*�Y��v��3�)e��|�����sNo��#�T�DIR�d#��:�������7xt|aT~�a[G�
��q#<�aAڔ�[͇�,TIzu��υw�����Z\�!������09֘3(;A�
��@uE~���c��)>����
u�5����Ϊu[r�i�p`IND�g�5ũ9{n{���}�<��p��v�VTo���۷@�w^"�M���Q�j��3��!I�#������$b�Q���;
by�1�Hu�a%mdRJ鴺��^){����G���2.��뮔����t!�8�@HV)���:
��~�=����o����$��ӉN��}�+������8n��o���gĳ�F?�E�e&��-�,�'�2H��3Rn]�)�KFN*���� �9��Q-,C����\1�����8��%������ɱ�J}�ۦ����:0���L��?g4.0�2>w?�J\��;�<=gp�.�h���[Y'�����_�^@"<דgǾpZ�{�����c������'�Li�D�(~b!�# ���x���o豓�Or:z�A���� �����Q���'��R;n�EOa?L�k��SԽYGG�-\�ѱ�C>^|��>�{i��t�H{�K��(�HIF7?u��Hu�~�)%�c�YG���+�yF��6@�;��W��7,9W	�z*>feP�jbG%�WᅂF��+
Iu���[eQh!]173��7#pq��g�o�e��a�#���m>CmbX��?��es# ��x����'��o}�"��H��r}�vX��-�+�QK>�P8�t�؉���(��������rd�Rː=�d��愭����F�-�q�vjA▎aTyQ(��G��U��/o�8<J�J��:��8j{U_������\s;\M�G�תg.��9���T�=�H�*�7��I�E1w�u��9s�4������#��D�bG��D=���2;s
:����TÛ��:/J*P��e��/�e8���ek�.���0 X2@���'�
z��w?ո��@�,�:	�F~v�6ҹ9���v/SL�A/&k���^j[@̀�(:��A�t���_���^g."���.k���/�߿w��`�e#�bh˯�U"�����3�d�8���x��e�ޮPAi�;9�
4���$hH�t�DY��'o���Gm��݇��C%>O���bYة���y�0�������ރ��j����H�8ɿ�f���B=bĳ5D�KT��L����V��a�qm>UJ�{��$4(��f�x>ԅް�S�j',�ڂ�'z�JD�/l��U��I��X&����s��	�g���9~�֚oL?�x"6�X��o8 #b����V��
d����t�$��&kf"!��X
���g�/>�˃��
����|���U��;���-nL��uX�����!7:�qb�S�I��r�=��w��]���Jk�B�'�RL1��N�Fb^� /��7,q0�gfWb��Q*�H��gC�OV�;��N7	��~�0�e���$����b�%1X?m�fy�
1�VH �|C�����/�Lb�2A�73X0���q�T�{s=�e�T�ҙ��41�˕mg�<L�;�%��}n:���Z�G=�H�2˴p�-�6�pJ�\��-b�1ߠ  
���
���X��D�r8=A�EHp2{?��*��1eT���4<N�e}��Ԣ0`�)O�s����	����'�"|>��;�σ��-��Ž|GF�L���/�=�N�o�x�o�k�f��B�M~&�����B�3A�t��0�wf3�-�0❐`��ܱ�Z�-UO���w&:��/�c����1�'i���� �\B� B�q��+��S4�}���(��	w��S�ԜV��{{�Հ'e v�I��{�~M%E�<�f\#Ov�������ȱd��σq�y��h�߃S���EK����9w	a�u'�r-�O�c"��	�tl�چ�|%{���X��q����a��m9A�44>W��o#����r�!ψjl&��5�$��r�K`��a�3�@�׋7�HgT齲yh�hM�N��I�0Zbߜ��k��f�\Li�@%��Z��H�˚��a0|�[��uk�%��0��	��g�
�;]�h�{T�>��-�T`�1x��F��<���5ZN�dT�O_��sm���>o����/���Z���=�\tjGz���d��g�y��s�sZ��bv���rbQ��۞Ԓ�	AF)�g�?��*q�Ҟ\���wXx-a��U18�FҔMB>�e-�to���+��(JC�����%���p�6���ؽ�jX����4Z��zU
(���G����\�0��snq������G�=�	'��)����YȊΕ��@-���R�lD�:��֐x���$���~ɝA�ҟ.���M���&���ȅ��L�n�8�bR�/�a'�E�1�p�M��W�'��m@��oP��}5@�C����/w3,{X�қ)��6��H�q���ܽ^@@�lhӋ`����Gӱg�pxH��/������{�Q�~�T��t��Y��=�c�n(�cw�yt(�|��'����`����S�@��&?�En�>��!B��x�).��~G�ۚ�SK���� �%;�OU5��[�H � ��X�}�[��n�5��6m��P	w7f���I��ȑ�'a5�YN�:z�� LQ�-@ ��~��{V�U��-�j2�a找��	Mq��aN-�߮[�37E����l�F[�]�kd�0�<�/�LB��b���Tq(��r��UWF�-"�!'��J�-�XMk�3g�/�P��6����_&���`}�P�s_����.�x`��!h�!�䢻��?���QN��mFoV�>��r
cE����H�|�'��W;���M�T\c�k��;B�������V��^��	.��Uއe,��F�Pt��(�h�� so�!�\z&��z��p 8p̤=���(� 93qo���^�֊��c#�w��%�=�a�1����t�M_dw��U��RԸ8��V�����Yl������m�{5S�9yc.���@�����G������Oz��3}�8/�ݪ �Y5�ډ����A]:߻�>*��9y�Ģ�9���R�9zo�cNv˵\
/�K3����Ď�u���^|*tUQ��x <��:�-�&x�|����Ybï,��9ɘ���᱃����J��6���t�+Gs�M��䄶BX&�R�pz���F����c�y�j �/أ����7��� )����Q>��)���齰a^|�i�ōHa/��[ўܛ��I�B�5�i.��qe���Vcg�!O�>���Ud��Q5?ﹸ�1b@J�'5�ϷC�LM+��.�d�5LD|��lg$u;������Ī%oʞ����+H~��8\�����ie�M�6��F����I[�6 ઊ�D�~wYM�+�>�r���A�Z�d-�^hܿ}��o����H�A�כ��}v70q
�Z��1ܣb���<�3:���2�M*�:O�M�?D��aH'�K�\�b��h �Y_4�5�?.lb�:d�^8���t��8\��ye�6�%����b�?� C{a��.@�){yUǵ�ޣg{�x������O��B��P��J�k|���8q�)1��}�d�D�t�E�%��f��/�W^?���.��Q�g�V��Kf�r^�`-KLY���|A��뇚�o"LzG23��ż��e�>�]����y=�q�;��ŷd�N Bg�.�	m`�����␣)�侏�571�����(l���}���[��9�]�J\�(���9!�.�^�1��h�7P�﵋*B<
�^�1E'����5���β�xPw(8GLDv���|z��M7�qo��%�(�N��e|9�20�P��O�0Z��loCr<�I,݈�z�K�V!�`0���K��#ݚ�]��^P���x!�Y�b:�fʪ��'�90��N�i�������J��!�3@*r���KQJ$�(�%�A�jr��o0H8Xq�	�jK�����K�	�t
7/n)i
:K���uT�f-��l���&4��i�L���oy���(Z��%��\��6y[ .�!%�B��&���~g���
����꺠�����������) �I��dWҡ�َ�p�x����g$ؖU�H��I�1���{��0����[��hR��m��P���ܠ���R�ĝ��ɋ��Tf�X�`G��|)VY�wwŢ���ʄ��q;�Ufh���#=�I���7��v�.,�_�v*�0\���{֦���
	`) V�iO*<a!�u��[{�ؙy��W�k�&�rTK�.A?Xp��lU1��W��9P= ��b6���^`
�{ݥp��/ȫ�j-����DR��p�2��N�>�]�{�M�4��t�7� "���FJ\����+�5��C�j\����D�� �}������� �&�vJU�e���j�a_m�Y�!Í]�P!�Õd��O?k�ņo�j_VB����,�Ǯ"��Yzر̢�o�TZ5�$v �+�&����~oj�4�{5%,���չ�̓_�/��%:�0	is��D�Cd&�3M�o��E�ǎ��kP����j�}��T:aڌk�ڇ�{��8��k���%4�����X���O�~�7L������|�轑-oPB9�20��N1�_���O�SqS)��@^4y�Jn��Q�`I
��z���i�÷۲!��	mF�zЛ9��&�.Y�zAú z�9�'i<�!��:Y�P��J*��-H5q:;��.o I����;�,g�u�u�����oX�-� E��K��1�~^~�H�vo��#0��� ���%{�嬠г'1��Â��N\�QL�����t|L+-�l�^0W�jQ���;���4�f��u�D��&^?�~�S�B���P�=���f�٢-����9W���5n��z����.� Z�a�$�������-��5*@�*�2`&N��󦔷/u�L.lB���'�ߓ(~�����1��Hta��!Η�S}r4�8Ѯ���m�@=-D�
y�Q]�"��/�e��+"h��//Z�
A�����l��<�v-?N�z�'�{���)n>�������n}_�@����B������T��F Q./����Ͷi<}�\RB����-�3{�����"��S�4>�.��_a۳<�,��֡���(,�A��,������ևr#Ie1�{���|�r�⛹qX��N����4�H��0�LR0��_Bs̫R�-����`?���9���K�\�%9��5�G�ˠXlxVHYEB    37e0     ba0������^(��6h]����r�������H�S{(�U�Luq;�W��Q���UZ�GI�V�@�0�F��O�ş�ؕ
�y��j�';���]Ht��+��J�<�����;ϐ��MͿ���g�,H!W޺��>�(2�5�>YT�Y�T
�*��)��%o�����d�@
�� ��~�a����9K)ڿ�y���RET�������cI"���4ڟ u��Ȥ�rO�#��ޥ"�^	��A��[Ie�ncM|�}�����1~GH��7E���X�V����;�u��:A)SB�{t����k�A�(�^�7(��T.E9d>P�������ʳ���Ĺ�#&B�zR�i���0�?���6j'_��q�ܟ��VaYr�'�4[�j�qm�C~ts��0/>��,�w�T�K7�S��Xõ��I6����sF@�� ���t̄�$F�6{�G������M�mw:r�QY��IvXTj]��R@3��z��)h��m�m�{������ۚ�Թ|��Fޛ&+H�nܼ�rxYX?W�� F��_�Y���F�E{?�y���.A��kF��>M�N%ܕ�)�l'\>�5Z�_�FF������ܞ������4i�@����s�V�pV*r��fT��3�6B2�� � ���9�S2������V� T��e`�1�FY2�p���AC]J�mRL�􁓎,�~d�����:���9DK�K'#2��	g���T�*��G�����I��'��f3k�+"��:�*Ҫ�t���ש����}.D��\��������m�0��;Ǣ�5�����;���Ϝ]Y3��Sz��7l����Zs(�������j�w"��X�^ݻ��|ƙ.8���KӨU�0(/g�Ė�~�;*��(�P�4���ٸK�`;#�G�����4&��42
�m��f�3�*�y!I�ؕ�bw�.�� �K��ׇA��u�p�B��#56Ν���l����9R�y�"�zh�C�S 0�8T�d͉�@�_ʅh��Y3Z=�0H9P8Eg�}�ƙ�?t��=������J������>+9�,|C��@`���WWU=0w@n��?��B�cn[x��d�	�ań)gH$L��)�9[P�w��y<��_6�oh�G�K,� ��2�eyv]+�L�M�s�ŧ��;'n���,`}�!�y�S�,[=��Z�Z/H�Գ�J�C�?� ������h���G�_�� 퀽sŦ5~���K�Ƹbm���?�]�rC!��� 
~�e��ΊqZnӠ�:��m���z��r� [^ۊ�������?s+�b�"��O�&�FrKѡP=K��t�|�R6�-*S�#�/ˏ~���@;x��H�iB����G�L��6��b�*z@0����kl�5B�"�7����i�8�	�� 2�N�'�j ����{vF���h,f�R�ot\��Fv�1^A!���Y,!D�W~O�g�waP ��˓6_�L4�@U_/�(C�w�1��e3�����8JWn�aX��m ��(EJ��!(�c3��6*�:�F�Ϣ���h����a{���)��Kr�b�#!z�0�;Q& m�7�)�$�{����>��5�ͫ�r�®�?�U�0����S��55A�K��)/��6E�UC������+IYL4o���q�:@;j��kR��@"��bW ��ʀ�z#d�x��!��P��"	�O�[��U(������k�	����~<QeԶ�'8���NerؚTF�jK�=K���V���ɒ�S�H�s�`d�U�g�=a���zB�� \ӌϓ�������\gC����dND�H5PВ:�K�۝HUjh���H��?���(�-���U �;�ջ������0宴H�����ȀQZJ��(`�q���)�YV�떾���R���������yv�)���%�O��f6�~�̓���D���ҏC��d�kM��'�`Yl��|9��N�D�UyNo�%�u�S�z����5����T[�r�?��~q!�J3 #|��!IU��J��Kv6�(�7*��:�dSM5�)F�gհ-�$�.�&����!�Ma�'��M!ҜKZ��g���+f��Qt��Y�%si��#i ����	?��ʷE� ���*�i8G�N��h��t���pm�j8�@t�呎׿}��~5���T��V^Z���-��w���C�ix�ܜm,ǿ���@�Ps';�č��I�'7ܔ}[��U��A��q�CP\dQ�6��5���1IH�Wϯ��6A�ó	]�.�p��L4#W�qB�kU�P-@���� \�K�쌫��x�$����G�kv��n�\���U��[cl���
�/�o�E�/�/��;��J�$�J3�
��p�#8��� ���Q�jU3���I��#q]����B�V/j��%ߝ�V1��)ǵ}�b�?˺��V�c�f�|g�����x+b�3��1�Cx�4�&ΈO�������	��!*3��vN��F�m�J��~���S@NS������C���7�Ǣ2�+��H]Z�A�f嫤(��W�[����T�=�i��S�@Ҥx,�AT椰����Y�,>RO7��}Eo� BB/�o�)	�9�;�KǍ%
O�j��L�XM�Ïz0�s~d3��?S��p���K��'���'�-`�o��tؤ�`O��〽�B�4W�_��8����9Ēw���3����E�MBM�k�1��4�Fs�G�;ݑ�̭�r�p���Z��
<�D�}��e��FK��q��(����u�X�/;ܗ�xg���x6����[69�7��n�5-��"ؽF+7�&vٸ�חF�ܨ�(|��x�8!_�VC��v�ܖ)0,G6ոʺ^�P��	�[�*W��쒞����It����p��y�����׭��wؓ�.����6