XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��P�x;�S�� �wN�2�5��t�,e��$iݎ�mn���u��OKc�9B �<�u�솽*`�_Ǧ��vѿ�.����i��<?xh��4�
�� �-�E��}�6k �7��'�,������S�AR����ѹC�\,�}��3�^�M<���:�k���<���6��^�;� �#��_nb	�i�&��_�'�[&y��b�|�0��;�97$�V�Q#�=�t�?lm_\p�Pc��A~m:E+Ԡ��:(n���V��ڬ�����\�w���I�ej�)� [sA��V����I�����%S���c�De>+��$�_~�E
���Y�y���4+&I7�>]� /�g@}���Z���2��3*��hI���#��g��q3�u�#b�bn�Q�x�1}�D���n�5+'�A �%j�|� ����S<Ȥ�Q����(*��H-���A�D��2�6|�؃D!\�#�q��A�}u��X
���2q[���w�k��f���������/ﴍl��ߒn
q�t�b](1X;������C�T��q=z��v�p�j���!�7D+�����30�p��"�6�Z��'1X�q�#� �.��iG�LgqS�AY�[R�5�;C�5
Suz�S�`�����C ��rhwbi�CO����T�ܜ����E�{Ǚ�×��4ٍ<]���X��R�^�����5�&_�R���/C�=�$5�8i��WV���2�T}��У��v��l��XlxVHYEB    2fbd     d20�Q�N�����}����B$j���S�b�J�|�^�0�[���N��#D�[Ә��E&W��k�S��q'��]-:��Z �b��������4s�
=̇�7�s��ç����"ǣL��L��K�1�����	�n:H2Y���ʍ"|a��6~�W��뙅:�6��%_0	�x�ϸ�*[Jd+g��uV��-2�y �������t-H�w�2��hڠ���ѻ���W&���l��뉚�S�nD<�����]�9���P�-aȓ��?��."u�ZY��kl��$�:� ���O��V����`EVhd�ؘ����6*���=7��;��5��}%굌���\����C������O���?:�c����U0�W���,�U�!
�j������PI(�V���aN�3���������'�� ^>i������H�J-�B!H��/$����.�0����kK>����ܼ��f|K�8	'�5��Y$q��mF]���*}�-�nث�sA� 7������f��ض6d�ܓA�d+�?6ژ~0�߂��������K�%�Òyw�E�K�[�!Eئ���{�t�B�G���������Q�NG�6�ڼ"t^m,zEWL�;!��g�y0��Tw�%;e��Z�R��x�s�{w�Jzs�]k�P�����WJB$o�b�L��Ǵ�pFm����ڨ�[��=Ny�
�J3)��d?_�!�&kS���U�_��]�8!���QM3�R�9ʮ�W��j`q�����n��+L�\�w�����~�t��X�+	F9h�U�J��0+�?�ȑ��SSA��!�u�}�<rW�#aP�MJ[���thziv$G�?���
�lmr� ���B�4����ߧ�e�T�@���Cح�r�q�+��.�0=�1�N[�п���vb�62%�R��s�LnJ�E��miuY�\%Ȉ��I�E.�GY�H�:����Ý��y`d�(��=����r���G7��y�
�a�X
���C�@ʅO<3�%xe����e�7M���צ�����`�v��辰&��O��}M�7SPE�V���/�r��X����y��}"�S=��ם�SD������޺�ĉ�UKv{�t@js���)}H�#�7������U��#U��C/h3"u���lzG��7�k�y�S��O��踘z��y�?�L6��/��Ԧ��3�`R�A�q�6$�%Ⱥ�3q��Ա����)Ȳw+.	"��z�/�8��WA�� ����T�x�2l�������ϛT��SXY�0����	0|jx_����n��U�VW���G
�Q���OY��x����(q�:wE�a�0v�6i��?j+oA;6���	�EG����*���+ӑ<j�@I ���mi�u���,$�f+����Җp���;w]��E��P��ӡ���~ٺ��Җ2%$��<�_��o�{3���\'��聨��)ag��̎��lo��M�v��MN����)��K����V}��JA'��R9"���t �)�}K�W�b���]⃝�-�k�_��6�yV�k��j���~	�������:�_D[��uY���E�beW�N6i����X��A�Vg�x�^��>Q�.jdH�a\�%ތ�����ł'�`�~y�&��A�S#���p�������U�?�6��*��ϧ��y)�ͤ�$�F���,[r�Մ��<Co+�aq����Q�����}#�<�Y:��w+-+gL�;��	?���1�6���eb�&�>D�.U�+�y�HF�Y������H�uU����N��.�z�Hw yD&��������[W�]�LK��E����^�F[<1Q�o���Ċ��w@.]�?�{�u9��+��h5����\s5��m�W��=��/g�Dms0�]M�ҜCTH�X_ב�,�=i����B���u�6p�y�`�
h���\
�@�ʂ���+���������J�7B�|��^�/f���s-z>������R��ٝW	%X���Bd�s���`��>��-�ȆDQ��5w�r1$PT���~p�t:O�����_�Z�${W��T�����5�`�����*����K��P�b�ǽL����J��6����8�;n��O6x'�����J����l�{$*vP)܂��	� ȲͰ��H���5�k��P-z��6��XEҵ�8F��k_wv��9���$�_��i�U����q<Cc���X	Q>�h�]�Q2��,�J^���:V! ��QA~.�n�k�DZ<gq��~|ŗ�7 ����6i(+��j�{�b�YW(T�1;�oA�d�DK,�?���3i��hun����/���ul�v��t�(��_�i�:W�k�9n��I��P�X_�m����lF�X��� 8Ōf�v��
o<"Y�����Y��(�0�~\�#D����J�� FF5�/s��l�켁��w< q�@Rc�YK��N�lF��O�\��q����%xcBQCWU%�>�uJ�M���k0�D�7r���9�L|�N���>d��5g�.Ӆ��޻�`2<1���L�y����'�� ]V46Ք�NV�~m"N�_�v ⁢�:G��UO�8�zڛE�@��'!"����@U�����#�u�zq�O;3=������<�����VD��0�����,T��`Q�T�\��ҵ?ǻ$���6��5�j`G�̬V-<K�wlP~PP���ʍ�͠=��=��T9��)�	����0^�;��_0��.���9�A@Ǐ'����i�o��w?0+o�>��>���;"tf��/�\�ryS�����S�Ux�N��k�c��=���9�0�5.¾i�+Hpx\��2�kl<L���;��1;h�#��jl7�㸒6����7���qt�^�ϸ�p%��o�:�ڣ!7/k�ʫh.�bgŦy�����ʞ�l��	=;Qi�KڎY��N�rd��q߮v�a"6��T?��1�x�1�4�j-SΞ_��a�v޿��wOj����+���aC	�;2K�Yu��V�-
4���w�}d}��g�Ο��<�Z?<���B�
���ڣ��y��5j�X�T-y����@�'Z}��'���(�����5�-��J|��UKf�￳��K����_u�oF�hv�����'�c�����~�4s�)
��rՒ�G�f��tQ��-ի�x߇5�����%������[O��0��ո�hs��w^ �������w���mV��G����F;����$s9��4�5s�$7���