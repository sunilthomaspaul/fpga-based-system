XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����!�F�����a%�0�n�q��12�TL�|�{L|ճ4D�?�,�Cx����yVȃL��-�r�(R�%S���qkY쇑��:��B�n�X}����g���(�]`�.L�N��ʣ۷@zD�%O.x����D+�	��Am��Q�&j|��L7���=�X9��\�O����<��|��Od|V�q�EZn�Wm�6в,e��p�i�m��A���T	6.�E�B�*ٰ:蔹\��`J�:)Wj��Lv�\z �V��T������K�C�M����*�(tH�V�a�(��Aq�� ��$t��S����}L��K�ޓ�[�}M\j��[����=r�f��ӥ���g0=��XB課����<8��I����op������V����#���s,N6��%���ɾWjr��! �A��3�$is�%�&=O���#p�u�{mo��� i�2;ej.EN������,0��cd0��5�D5��G63b�u���1s�����Xp�$ �?`;�?Զ��v� ?�
��J`���J��}ERh���W��������/Y��%��n<�� 
_��O~�PT:�B�xL�����ʤR��-��p>aJZ��/g�ێ�`��(@�r u����!�l�oZ5VpK_(��HÏq۸!C�z�WH���?L	����]��p4��"#f��'�wlMO�[ǋw�:�!&*C
��p:mK�h��D`z�q#��d��¿�k�5��9dXlxVHYEB    5658    14e0�<���°��~��5>c�P>�/ڥ�R�^�k"AP��a�B�k�]ya>�!l�$�H��i`N���R%�#�|d��_Id��W$���~&�#d�&����k������\����gd+�	����	uPu�Lhh�t�������F�ǝn4�9�9��,p ���ށO$�w	�݉��J�'c:F�Ҙ��=�H�r�ž�]f$ƪ��6Z�X=��͉��X�R�\9�(�:�7�
�{�u��HUP�Th\�����Q�Kz�{J3�To�rv��  ����!%�9�]��m��8���7��ح��9&t�^�(Or�CL;�el�tB���<D��M�w%ę��R���3	^�N�(>s��m*��*�g%��P���E���A>h6��(!�V։K)���	����XrJ��(���Bڝ'y����=��*k��!�t��yMg��'�4�+ƻdT=���F���ʅmj@�c��1U	�9�ۆ>	�S��UkD�.��r�`�Ӧo�O�q7��8�h+���'�$!HV����qR�2kϒ(��+�tP�d1�AS��l���:¢�Ά�;��S�Y�o �
�@�nFʸ�feú|k;��� �<��������H��bĮK)>������6�m�-���k�;���j��.s�ܽ� ��ѐ�s쯙q��;Q��&�7I�VKV`���Z�%N�x�q�����,�ӣ�(0��+�+\��6�?y�^��0a{�!	�$�wO��NUڃ�݅H1�]3�3\���/An�e���'�k���0�b��3uc��4�5�F.��ϰk��c�|�N줇[��@n�Ze�r��*<����y����٩A��5} "�a1qǍ�B�-�N����(�{�ʦhw�
��z�5���_V,�%b&������b�2b^X&)b:��4h�5���;h����\��},��d/+}�&`Ɍ�~EK;`�Tkf/���E�N�>�z5���}��Ň6��o@���� �ʱ'��,�H�h?w"n���R�@�yA�	�b��"�@�_xg���*��c�����7\��Y?răUu�kzn�Hr|G�U��	��@覍���͒_��O�Z,���Z8cz{F�<�)[Зa:���$�U�9M� k�8��@K�^��̽Z&� Y��'�JdAR��3r�z��{`����'?��T��!f�݌B}�B����9v"Z;�@&��D�a���⨔���QgIV;�D�.k}�_�-/�f>��:���-K���I�4t���2������윀(�,*�do�h�#v�01�b�Y����!�hw�3O4�I`�Q�C'sEB�H����sJ�N���{
R����#.z���Fz|�e�M٦��4%���s����X���1���B�+��O�	�D������_�*��q��i�t_�H���	�.6+M����%��+X�S����0�&�dP�B��<q��su�u�MA�t����P���#L�(_�G(�qtې��^n��)&���b�@J�y�������M�����kܙ-R�)�Z�ŵ�{�/{�kuj�����qOk�y���/�mĥ��g�$�q��7�U�S9�n�+0��Yǉz繎����|���_��O�D��P����ߢi{��iyT�ӟ�R�� �,�mp\C�T�������y�ͅ�`� �i�rC��A�����3�B�s�O��9f����q����z-�Ux��F��^BԶ��D{��hpCV�t��B"�����m�j���-i*��M�B5�2�~��-������*���K� �Kx�j�ٚ�RL��,Գڃ��[%��U��s֪�����>��9�-:d�B���;:��7ZH`1����ٱW�{L��Q�|Ʒ#�Ҵ����W�yMy����^�
����VvJ��}ŖFq��Ur'�cʗ��!�ӾT?G�hI�%q�v30���+�4;#1	�)"�����{3�(���K�H�����G�#��͌�hӵ����s5ڞ?�%̛ �Y��X�V&���U��tp�췘�9~z�1|��0[�Q�A��Z| �����m��6�³&R�uޣ_��3FQ�G�s����)��n��,��mt��K�T���D�mB�~RI����u��&��C�G�Υ ��\I�o��D��-�@h�lN��hz�-S1��VO��jr]K�9�D� ��M���G��hC�H�n���&�	�S! �	s���`̯�:'��@3���f&�Qq��[#/��V���VS�ZbQ��b�����f`9��PO[��c����	�� ��O�#�G�Fx��\��˔�S؍U�=^� �zľ�>�&����"�������KP<����U񙋳�Dc��[���kI��_��K*ޣɫn�D:3!�����&�7C�JG[;��Qq�+��}���s�ڸΣ@�uyl�h�Ao6�AҮ۔��A�?�IN�D��Ԩ���鉤~]����@��3iwb6���~�����۽Q��0��q y���vq��.�H�c��rV�w�G���'1^�E�ֈk|�7A��ɇ�BkH�
�q�%W m*e�p�X �IYY�|��c��{�SvC�X �gr�7�����S�JJ�ܧH�_��V����m��O����
7=X�{,�m��:@=;5�@whT�V��3�U'�ZΉGBRۧ-r�7GՎ�����t]H�֖o���c;�}��Ke
cMS�7��Z�$u�"m�./pw�*VUԳ$�dV�e��0���94�lh����@�Щtԯn�TDrم�\q,;ʴ�HE��[��-t�>�5+���wm"�?bmS7E�Ԍ�p������Y�/:�]�Pe[�q�5eX@i���jaB���*7��҅���w��ĩ���W8p{�?���ő����ǽ$Z+�6��=Q�˞u�Of�y�]%i���\ux|�YV.�o\�?FR��f� )բiۤ��9r�}J������`$N8'�f��6BF�P�Q�7�u����[{�y��#�B[}YF�8����q�ze�&�y��l9U�{�j1��/�{[7�惕�}19%�b�	)���]���,:�Ӭ6X���I�K��q�O_/
���k��&����W͙.�i77���(��q@ =�?���e�ob9�dO��4���D�ۇ�O��!�2z����㙐o�+̑���O_AEL���{�
���V+�Y���Y���aj�9�N+�ކ�^���⵴��l��է��0�㢹ˍIꨖ�I\i�����e�W5��=B�a�oI:�Q?��N^+�/,���2*?7��
�!�%���if��>t�@���w�B�\��h�FA�2�x�]<sgZL��/9C�6���Ƈqe�=�
uj��h0i2�+x4=L�2Y�$�`�Kf�3s;)�BH*d72@������,�BD����7����O���O���\th���}��A; �Fcg��Tš�����鰜)��6'J�q/�`4�˯����^Hh$"�T=,�9M�i�PĢ��s�RE��O�C�3d�~uɪت��46�q����*T|���0#S������o�����-��I
�~D7�)2Iw�p8�Gd�e%��IRCc&b`8;4Rex%ѓs�ĥ�����g���<#�����g���;�3s!�=��=���ճ1��v��9����N��l=��W�c(#��c'A �?���?>��iL��ϰR��~n���B�Dv��xD��W� O�9-� F�s]ǰ�'ST���4ְ�	02)d�N7n�/���-`���B��<&j�i�lK��m+����+㹻�P��Ҳ��?tL��8�^G�3���[Y����"���ݓT���R�@�Ĭg�r_N��\�,4C��.5�Z�{{�X��� ��"#��5�z�]�谜�����s�8B��U�ؾ����,��+T��4j
S���TU��K�zq7͂M�	FS�"�����O{k+��ni���i��!����{\ȴH�y��,�X��wB;F>�n=p��n�7 �(s�+��TƮ����%�qx<k���B��Mz��$n�&�)ှfB�����USn�.����)#�p#�J�2�H1��t��~��%֔�:�oy���O�d�m�lFr�?"�����}_�;�@X�- �k��_���VO�B���|�K���nQ�靽��d���6�Wvd_��q�&��m�Z�$Q���u��*t�ERqc�>�ȵ��=��2W<U��ۧ٣
�N��Sh-c�æ�HQ�y[�������<�K��ۿp��J��½�]���~�	�	�M����JB�)hX �؂�\pci�r���p髮`3H�-��5P0W���Km�l6�!v
>�F���u��b��=xҘ�_(��T�ܯ�����P^Z�v��6p�u�hGVL�2��P;�*�T}K ��e1�۔�r/�B�Yd�ͫ��*sx(T���7.�+��I
� ��-�cu���/��H~��c�����p�I{}��+���Nj[|�$�3Si�C����hw6�O�kز;s�
���8���5��v��$�]?��v�d(W2�Џ!�1F�y��(k�c��T�"4���	r����M8�kt��/<?��;�F镬SaF?G�`6�����?���Գ��B%yL�lFe(�4��0���R���Ы��2���8�i�E��)�����~�V�#Ox�������>
1�W���*�J����;G���#f�D����v7� �$H��I;G_����L���|c_�;��ĉv�����^`l
�y�(� ~�ЕoLKT��v�e�vrgE��̩C.�dt_
�ԝQ[��2+�:|~WVU��ۖv�����2e=�����D��\���~DEV}���_ 	]9X��%�x3��^!^%�	�����0�fe�0�}I�&��$�%�q2�8���#�x�o���ز'��BX�W�O��ك-B6`�W{{��Y,�l���U�V'�ʥ�x�7�׌�/��׿���iRE3)/@ߌ]���,K��Z��
�6Qk�
ض�vm�p�*�}zx�+����E�d��%��@�����qF�d���̺K��;���]8�� �����7���h��M��]J��p�.��0�