XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����
Ce7ʖ:���b�XU�0������R�"����>u�� g+�H7)��".NE�q�g����Cǐ��#��OWo;4X��_�k�����?�c} �̠Mx��2}�݈{������Yݶ_����}�) S����G������{�/5ո�&8�CU�mB���g�__����yO�D�h�H�x 1=3bX�H��8[�& w:�d���v@��Đ�ѭG�˘�V��Qn% �$��rE9��'��PP510�됕֔�N�jb]�<�cz��R҈���D-iC4f��E,K_ ��gy����0Nyv6�ڟ�tS}�7��-�Kg������\o�Z�����Ӳn�Ӯ��
%��4A�����Ys�;����֏*bL�h��5�{Gɾ��7q1��	�&��J_��.��_�S:��S��9�P����
� ��|+�n�DLR��T�����3=���W�ŨY�i�p [eq��ʾ��qL��RXL�/4y��Sk��k�WYB~�ɞ㍛�E���o����Tɗ�1���h�/Y�V�2;�=�MT��Ǝ���g�y��M�k7^K��7?�t��s[��:�[k%M���ئ
�:?Qi.��>Qwwǧc-���O�Eդ2������oL���xęf��S�I�LX�y��'kD ����2�^�w��vaC`{q�P|ņ�egv��Am��d�.2�i�5�N�	�i9�w�V x�#|)6�:��c(�ѯ�;�v[:�]��Xͳup��XlxVHYEB    4564    12709٩0
Ԓm�d:-Je���m	.�Gߍ���rb���	)ԉꎋ4(��ӕd|%��ЬW���3C����xd��F�P0qGJ4�`'�h�Q�Nk��Λ�+o�ErM���᱾]]�LY�?N�9ɻ�w���J喪.��D.U��w͛�l����P~r�s��>��[�f򫻣�S03�۟���áh�RD6��I1��`�ã�w�����"jZ��/��j��
�e�yC�_�;(��Y{���(�����|D66Zd�pg��F=^��v�2��(�t��֐���z��վQ,=�뻂�m��ʶ��}m88$`��(�o��b�R?��_Ƴ�&cC�����~�l��o���4���K=��`�ǆп��}����uӋ�=�$fV#��2��EUx�.9�Z��c�֒���K�8
|^�
��H+�Y��EHW����s�Ι�rbhn*FD��+�ڎX�堩,�g���<ɳ����^mK?��n�Uz��r��>6kV�f0l�uf
=d�26�Ò��oq�%���1B���Lx�|�����"�^������w]�ͬ�� ��j�1o�w��2��t���Et@c���1���ތ��1f�����P���1�ǝ�5�6&x�iP��K��٥�
4^��6J����E@��Y3+qo��9��������s���4��ty��ѥ|l�t6]Z�^�7Q�����pe���<
L!hA�1�9n�=^ى�{�8㞖�1-�r�����ryT�t��,�Һo'�/{�l�KK�d!���F�D� n���k !����t1����e����s~<I��<�V�J4W�Q3��e�+�gQ�]Y�^���%����{4���Ykq��6ġ�!%�S�U�aQ�E��[Eu�q#;�O�0�n��4��Gϫ5:Ѭ]m��ʵ�ռ�"��9�#�Z{�&������B�'�D��
1�Hpٜ8���B��t�2.1O
��\�qT3��4
PZʥ\mtP��X{�#��PU8��I[�+�^����w��u%�t8նW����������Ϸ�age��+R$j�z0���� �|Q-���(��|WoƤD��7��~��1�9��^���pK2~I8dhܩ�8g��i��ᨒQ�)b�/J38��={k��$�)�}�����z�b� �	����w�dw�]��"B��c�ܿ�jZ"�E���l"�]���z��j�&�/J�����-��.G/�Q��5�SEej���f����oz`ޡ�EIzs�ٕ5yRd-�'�(������&��>?�����F:�l]V�� {4��t��2����.]�!"Pd# F{�-A�h��.�bw���)F��*��ѡ[�{%�L�;���T��(<��&b�H���#o89-9n����&��û�[Y^#c�Y!�������F.����,Ui2��H��܀��a���'��Kg���?��ʀ4Q��W;ʠu�_Z�<��Qķե	t�p8�P����c�;8�Y���/���3
-DlR�ۨ��_�G���.uS>:��b����5�6Z�R�\WɳQ6�:� ,o�~E�v�S��(L��x�.V��q��~/G]MU��X%����m\�����e�������	����������)+T�y�0\�(�H`T���aYl�6���$�`�5�����:l#��( ���o�K�+��2�U�y$ߑc`!�ژ0~=K*�$�5u�����\�%gW�{����͡�fgC��� �1ה@(t��T{w�l"�	@�ֿ��j�����9Js��W*��<��p��Rd���y#o���$�L��mH9u�T6�߫�U��z����q7o쥲 Cbm�M����'D]���1pŉr���m߶��PPtCV�U����oHJ�@���Y	�d�wX����c󞩺t��8�J~b�;�&�ȫwv��O/+�_Χwx����q0Z�r���D�u���+�8�J��q����qN�5v�[���=.�m��ut@��u���`���o۫��)�d^�����q����:x��s�}VK�N�	«�C.��'���K�	(*�h�$�/Z	wr�+��8� �E��<C��w^�]�t�-�k�ҍA�C�˃:��N	}|n0��B��0��QB�0�q�m3��xV��Q�qr��f������܇ן�;�g��5���B	�G�Z7LfC��ur�&űr����Y^�m,�r�1͡)K���%T�0�������[=r>���^-s�W�48�fp�b�����K�xP�IG���O^��K>��ǖ�O`.x�P�z����NI�207��:cYq{�����2?P��Z��ee�қ�|��sd��L;���
/#n�q(<�Z����g��.��I�T��E���1B���n9L��*`Gx���N>D�cz,#��Y+#�e����oQE��Q�Nʧ~&�:(��_C�<}-�<*M@���6���w�����#BП�m��}���/�O�Y^S�������ۥ�=_:>6��&���=�>T�	v�
�h��B�˚��g������X	�j��@,#)��T��WY��l(�՛���2��K������<�;ۑ���Η]���4�&E:��R&���&�B��ϚZ�pih�u�D���x��}�v.�ل|�-_,�|��ֵ+�IɹIM��@9[���x����ۗ/j��QĦ�zm���@Q���1t�n!�tk�h2яL�#�D�1�Bǔ�F/Hy�Ś��	��s�� T*�3j���Yt��H[���q�!�3�N˨G�U��5��}\1$��x�P����sv�Z֓	�(�	wx�0�uYOY;�.���sD�1�5j�]�.�=��9��eZ?J͈W��T�H;�D�U���/�Ҁ�<�p�yZ|��1��d����6��M��b�&��H��{��I�N;�m�+[7�b���	5�����z덌�2A�g�#��mCV�R�"���n��1�e�/B���Tu���P���G�Wcy��1sh�����ҷ7A����3#L� |����K�.~�?�yt{���$��R=�ͮ����#��7�dA%��w��2dT��q6\�&�͋��<|�qQ��}wٰ��ߠ�]ͩ�p�*��4�0�υXV&.̪�	�.K�	^��ʹ�R0�ep�= ��X'n����}L?0�f	Z���&�K+�&�3
��[+A���PV���iG2V�� ��NY�P��6�E��<U���Qg��Xq��׍�:�u�%���@xz�l�>)��Г	ku��ᶧ��kD1���F¶*�pR�a�q�EH� Ӽ2�j�f��z7�߄_���\0k�ъ�;�%���FZ�:�_4tw� �_�;�X���:��ܠ��r\a�N؅��b���赙��0n#ʑ��'��&.��'�<N�����~Br�$ �.�bC�N�^q�V�T�g��.`�
��ȴ$�J�C�`��m�:���_��^臰�]�쓈��
���a��ps�
lխ3O=�=�0���3��8�����\+��.�Fn!�)#^�������ɡ�{�+��m[��a�1���y5Ad&�O|��tt�S]�|�����Yz��p����N��g<xބ��l�ݯ ����{�8?�7
��K��m��I��W�i�� �"� 	E(Nk����D�
�r&BO�Ql�f]G���~K<p8��5�_�%s~���|�� ����fr=8=��#"
���C��j�9���'o%�
*�U��7@�	�����ٻ�9m���P9��_ A�����8V
�[$����|����^�\g�6յP�^����0�2�/��y�6�Tõz5����2OұX�{���?�]��[	�����.L����L�I���RS�h@unY�͉�e���}\T�@T=�0��yB���DS�B�����%�7���P�Վi�>T�7���P�j��~ʧ4����^�4�5�ʏ/h��8s����\(���}����b��|�*�<�y=H�^&9K����pS��G()��
J_���FӶ�ά/'&#捶��Y�!��;m�?,�|�~s�A��� ��b�B���K�D�����������[v��2�I�l(���A#4��p�B��F�c�RTAS��޲���?^��_	J�S%
d��(���JT�7�a@�Uk�-����f�Jv��n��<Sm�_Md���:w�p��G � J,���ťO�
�1�@���,R��56 v�yn�9��ts�a�5��p�����܁�����a�N��Z�$Ù���|�3��T��{;$���QA	^>u��T8?���[�[���O�9F�����4�iz������ؕ�Eù~ʺ|H�Q`�V�*�z庽sf1�(h�7��P�� ."�>�����g�\���s�����E��U�e���Ғ�y8�OCG0~2~�/I�x�Jϑ
��e����m�A{�	U��4d���\w��燶�"4E���$���I�kN��Ml���b���p�D���!��7B����d�����ajc#2��'������w'b���n������e�'���#=[��ʨ0m�)�9��LGE���;(��_���(na���!�I/%�L��Hß��