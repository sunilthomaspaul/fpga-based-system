XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��9�X�S�UƘ��ŋ�<��p� ���� ��C0�YgH��ܯ���l��C<��SI�:A����x�g�)m?]up�[: ��K����d+א��_Fڿ6rI�[� ��N�?#��X��9asa�:H�L5W���$0㔛3DȾޅhP�"+͒
��&2��7B���)��R�k��o[(���S2���]<�9��R��r'{%��vd���d0s�/���ucP`�a1���1��r��93A.��.��tӻq�q�,�(.��[��F���b�4	��r��*�a�¯2&��np�6{�)�0���{�}8�T2�x��fMR�F�����s;��x���{W��*D)��ψq���W8���@{�Ǉ�^@l�D"tQ�Q�Z_H����)_����'8�{����`�f��G�!�c:���ҏ���&z�,�蚓Q��8�"��(&t�W��Ο�g������A�nrF�m�M#�/O�K �x�^��LK͔��u9�M50|#�<��A���APKt��#��gR>v�A畄����
���.?�"�
�eru�=�9��陗��3�O���'�����V��s�`(���ʡ�6�\�@R��c��yřa+R��0�b�mur�(�"ܩ�������R�<m��.��d���p�����l���'�� 0l�����O�c�E���m&���=�_H�1,+
6(��J;$��3�[��c:��S�I&������I��~X�ΐ��Ϸ�-XlxVHYEB    4548    10a0��Y#o�ƨ�-�hr�~D>����^>(��hq�~S��0�"p;��o��g7��k>��>�h�.m����1�D����I<�S�^d}�5�J �o�iAf�X��G���|���n�ZW�����p�
3�j��jS��H�"d�4��T�Q�����:�̣��u��R��]ឮjb�oc�Cg��7�pN��fxp}v����s�PXq+��0�Dr;��/�7�r t�,�_w�͖#��M�jT- ��f9�h,/����d�	�-ݾ玉��;�Z:l�L�����������f��m�~��De�+Ǆ�dѺ���E��}�O���.�0�����ЬCN�H75SG�,�Pɹ�6x�X1؟�7X&��ޮ��\�R��+M��g俣F��|vp���C�(�æ�­|��?��S�ʗ����j�IPL�D`,x�TkM��[��+��(�M�����>��j{���8h�B
��1���d{=�MrW�>��)��	줂�G`�J���Ծ*��p����$�~�<����8b��1����Ƽ�Z:��X#L��W�P�+�N�M2��0)�t5���5@�p�I�q�^�ܥ��������
.���	\L���3)�@>	_N\�z�h��y5���T�����]K�8����UGW�##(o�� �#����fUd�(���v�=o�Vڱg��Fv����q�y���D�(��;Gad�d$5qH�<߆(C(��G-���
~�<��Ze�ة�%چ��)��;4wX�Y��`ݽ�|}Kz�a��S�%4��6���-t�ҳ��L3'���,��I ����;�W9u����E�Q�0��W�?�f�4*��.� ��Ǥυ!+����)x�t��H'U���n!��B�Y���s���e,�yf�NѠ������Ą���~r�v����U�?7e��W��d�_���S0�}*�Ƃ�_��I�14�;�>R����p�z�7��W�s��4�V�o�
�:��X��C�w�U��0T�ڮ�U[�����oΐJ$�I~�{�_e��;��9[�+6'e�#˄%T{R�!�_c����/����ݥ��fڑ^5��rT������	���)�oí�\O���Β��I$g���-Q㵲��?�	����z�['@�E�$�Aq��6_m�b�2��������Y4��`��&�� � �R��Tf������V��{��>DK�Pxx��O�����G i�K�]�X�W��ح���T�,u����g�����1�7�D��Rx�mi"���w�c�F�u0�Y�������"C���	�~qD�^f1!]���Ȫ2^� [�����*�Y�;��P��m�Q��u\�W�/�����}(A�=�������v��g/HzM��*hC���7J�C7���� Y1�hn$B�)�8���M*�zl@�����/H�ϣBs���m�B&A�_ú
	�o�ui�	�o��ؘa}��Ć.�}��=�a�>��@\p<�;C�Si�d����0�3�;��â��=W(��I}/B�h��;��q���BG��3=�������Һ�d��+�v=��X{H��ڀ���{F,�Sc�v�Ϲ�������ĩJZc��2�9;;�e�CdR.�����o�¦{��%N��/�H��6���\��I���%3 ��
{yq�5l$�P�)m���BO*h��Ӆ��/�9��-ᗚ���K���$Ng��?;�4Y~r���3�jq�R@P�P`����7�:c+�('7��.0��֛����!D�?�a�^wK��{m�M���b�a��W�$�;���,ූB$���6����i�Y�o�⺊�x�{�sV&h��pq��^o�Ȏ���xC���;�/mw�:R�����w��F��B��mσ!f�~�CɘES��0���:��8TZ�����j'�Ǉ� 	�v$b@�잌��k��1�X鼊'���2�p0�mFq#e�l7�'�mie��D�'@@|����	����R�-(��	;����+-���R�+ƒ�8�)��ޘjE�L9Z��ҍ�a��sc��ς����q�.��L#� �j�����=�s6�O�x�,W�H��2M�I�׆ֳvRآBj�����+j4�s`U��+��y��\���l�Hj^���%8_� �At�n�3����F�`��� ��{%#�|ߍ�S\���Xz�N���&�|�}�����H��HR&!�Յ�/��>��+rSف����"Lh"��������!�JS.ìS	׮�������T4��$��z�D��������$wn�ʋ��_5�z�ո^���å��W��۶�4"Dt�e�H�d$xf�����pA��{��~��C�!ju��Kh���,:��|w��	�6 ���_k@��Qy�o:���`�)g���Po����xI@��`��i>�x��	\�35�1�Q*<�Ԛ��C��	����j'��{``nI�}���R�+�����g;�Vs����{̉�����]���������c��|jMC-��qdEѽ��T�&��Z��`���D\���������d.2��]� ��Z�� ����A���h����~��}��s��a?�5[�^k��>��jI��y�f����6�a�ro���o�]�ͣ��l�0�! �[��������!� C�;@��(?F?��x�3��fԢ�F�4E5�|��9#�� Jv�@��6��S���\)N:�������{��FD��H���/#��7i}úBYUq������5{��Yd.�<�yg�Z��c!��}��O�@�X׮#���_�� ���#�X��T�����H~�@N��	�{�w���RWͿ�ֹS���Q��;���|����2N|�y�`�����'b�3Eq(բ�s/-�FA�VL�K�;I��&)Ԟ�ѷ�E�z��d�hm�4�ǴzY�v��-�@���ź�\Vm(x��w�@/�NWm7I�^?<�T�񩑓�	��ª윊�p�Fo�Gm�=���@���+C����Y�"�t��rG{��z7x�㡖���̛�oIc`P���o35p�ć� {ߞ�����ϕ
�(h�^�}U�Y��T�$����3���� PG{&��|�, �4����	O�y<�S�0p,��qLy%?SPF�C65�0T0&@=�����w�e�r�@�������ϯ,�=[�3�nX��r�?�D�/|�6��T�c��AG�݆=g�/��DO�x |����El=,2rqI�N虮���g��u]{�l�ϯ3`�	��ià��j$oW'ee�R����HW�n��)�.\��RNJ<�# 3w�+ե��G�n����3-���fW!��_�x�f�l� ��j]ObbR5)�=kCc���.����D��,x�?ζ�>�!G }|�rq;q4G������,�ɭ�Vj���D��7��\�&58	J�d�8=�x���)$P�/R)����T�Q����e���и��o�Y��x�LS����.���ŉ��Ș~��7�MN���ű2ӃsLhA���5�e�ER��C�'��`Phȹ��bt��=&�"���"_�K��o�1��`5����}�)ы=o#W�����v�� ���^4I{������Bw���sOn�8�j�'De����w�[>@\���=�C�����F~�4��X#Y�O��w�96�G1��<zѻ�<�;��O*��5N��5�5^�NU�i$��M�e�^H��Ŏٸ,bբ�ۗ;��<�������eDhq�����ca 瀖?�Q���.�	�w^Ȧ��ܭ���OUG!6�ʤ?z�+Q�]�7rBń&�dW�XD� /G6�_�G�pq��RS�[	�(2�D�k��m�����,2�����$w���rS���쬓>��v�8	dG�;Ӎ�ve��ט/�&�X��R�ظ���� ��	��f:Ca`�p�2K���56�	��9�ɸi��T���{�5'�*�aa���i_E�m:#g{�^?���G��O�dz��y]���o
�\����E�ds�s���t���*��4�H{����oks�#b|���nX��<�ܖ[c�S��]�]Ѥ_�^ZaBB���m������