XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����w������P����/��2߁p`rL�}�`�԰HR"=w�Y������a�Nl���{�k:�O�:���Qh����đ7�뢠�१t�>㥛� ��­�@q���U���F�8mz�k]n�5��'���3���C���Aً��<��&��ݺ�OM9��dX։�JW�L������CiT�$8=s�?���}j�u8���Ϛ^
��:��4��@jv�S� &�|�~�*\���:�ݪr�uw=���Ҩث����>Ľ ��Wv�Oy��_d���*��i5�/ \SG���W4���1�>!���}�%�U�|FO ���J��E�y
\С�������~��bd7<�Ղ���T�Z)��\�EV���@'R��3�Q���\��9N��v�����^�Us�ϧ:"�AB 9텓�z�Zʇ-G�s�+&�'�b��]�p�������DUJ�&¿rZq�>$	��H�G	U��&W:�r������������I���3�n���{iW�]i����� �WG!��/�m�_��%R�R=Uz��K���Yy��!i���JWG��3MW�f��R��?��������HH,h��8�+i�~�	����{"���7p��-Xz9���ڤ��m<>D.����$� �^��c�Z��(Ll|�D�B�u�:���:K����-�U�D�6Z?T��F���ɟ�y�Q4[U�9��Z8��=H �� T���(��$o�\d�*8�_�����ts�s��XlxVHYEB    1111     710���8��!`�^4I��5����&5Fw�;q`��}�8�gf�"�g�8�c���|::�V'~�� ���a�g�u�-��u}tVQs|Ǎ_�5+���o��@YY�x��"�"����&'���z^�P�]�$֢�H�$�kp0]�g�\c�6�3�,e��%c��u�T�{c�VJ#w����L�,c����_�v$�4�8Rҳ�=���!���cH�s���9�W�(I��)�cx!��lw���w�*�J"Y��: ud�F��9����l��u�I8���1�/m(�n��l�ոjr�V`��u\�ԣ=wE-�P��3�2(�@���cqu1����J�a ,Aƽ��	��a[Ve�!մ�Oh�����_������?M��֟Y7.������փl�%Ĥ�6�!�E��z��:N���%V�H	ǅ�����@�&�jnJ�yK��r�o��Ð_y��u���}���Ij���WTc IT�)���J��arn{��#�P2$�гy}������T��Z�VƓ�=�{ �Zf0��.c*�� ~$�"B���/]���w��B�I�D�G�7�8�O�,����$@pԙ/���ԩq�n1,�!�>	���k����1xG�Z�޻���9�����$��}��-<��)��70s�ՀpX��8��e����s���|]K�܀�,�!Vj��#�YYh${x�޵hpqc"\���KC2��&D�S	`�v�����-��]�ك6�_��{A�Ӷx��dtJC[�VtΔ�Ԓ���_]��z7x�g^&�xP	���G/ޥǿK�r���┛��=#˚�C�%b�z]�o�&%q��؊���D����ܲ��\8����4���5�!c��m��*����K۳3P�q�Yv�!uT��q��=��3��y$�I��^������m�}
�ˊͻ�����J�K��kH�痺D��g_���6$�q��~^�v�'�~�]��&�u�3פ�W?f��K{������A\�<�Hp��]j<�;8��rr�[�1��� �	��>'go�� �u�p�5k�Y� o8R������0]25fI��X�a!4���u>:���9x���?��Q:����..�[+��R�i���HS5TOK5�a&z9�5`���w���l ��G|d�� 3�Р�C��/��ёd������"t�`�\�ƜpK뢹�n�H�,��߀NL�[�N��l^z�,ϑ�Iܑ�!7��)��5�H��e�\u.?O�˛�&�P��dl?���n�ϖn���&k+��t�Y��	d�I�9�{&�
1�����k����b���$+���LĒ����ltgo���}�0^S�"�1ʻ�P������ᾎ�-o�|%ֺ��Ɣ8g�ŭ�lVV����\;2��)�=@Y�����5V����V�8�*;� $d���x��2%�eS>K�7�)�:=���;�qE(�>]��x���k�0�jDt:���f�֜}���Y�[�_^��LG𬊻?��z�1B%[�HFcR_n
�4�	Ɏ�W�ov�	�?<����S�K'�f��r�堔�DW@0�ڟG�o"t�XA�_,�q$?࣬�8ju����1��>?���17V-���	��ׇb�[�W��ԅظ�t��G>����G�C�W��:^r�C84�:�T��S�%��Z=�g[�p��igtթ�: @�u�բ/�.O�V��(��q4���M�cbz�8\$5,H�ujba�%�Exc�2m��-
��ȟ#��u�$���oM�o<~]�|��"�0<�r,�.��f4��_