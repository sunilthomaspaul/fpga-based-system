XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��R���^cYe��8���U<H��N���9_>�X�B:O�����P'8%J��[F�Y��I����� �Y��dTW��=+�d�oV��cPz�*��PwT��l|������^'rt�"2LS�8�	��_X�!9���g��ko�ֲ�i�M[�V��y�C�q#�B��������r��x��KQ�b}U^��*�d*��B7	)���M��@i�s��ˊ���k	]��ɷ����N���_��"�Xj3��%�OzH��wL�U��b�x���'�?�r�����k6�����M�L{$�!T �!n.�5,��Q�M�j���TZ��G�����D%��q:@���^�H�74�Zy��a��c�ϝ�<���"?<�r)������ǥ\�5�Ds��5���Y�W�����A�2�ʣ����M�n2�{k��f띧�I�$�u����Ї�� ��J�p|��^��NDN�ae5�'� �>�9���6dP�A��"�y=S�o	����(��ʑ)�wmY���e��U̵���(��7��S}����˷<~H����+K���Z��.�t���ټ��#�$�C�}�r�8x�3oxA�1\ɸC�L-�I��\�Z��\� �Ç�ˋ�OH�r������q9�hbq;�ӰG�2�ȡ����#n�Z������O��3G����8�嶔����V�� �KQ)��&Հ2v����7c��L:6!xe	��}�{Qw�=��B*�KyP�
eXlxVHYEB    bd1a    1920:9��Ġr�R�!����W�,� s��[t	���E��^�TP}4����պ�s�_���s�P�ESfdұ�p�|��Z�7���a�^�'��-����\c�3FI�EB��D:2i��k�)�PPa@�KZ��mK��pD/xw�j!�}h�������S׃�ۏ���	��3�-l�ը$e�~�e��>G U���̍� �8��ā%�7��\����!I�〫Ih#?�(�!<'b��g;oTUvt��J����� ;���Oe���{d��H��a��Q��׾oB�,u3��B4��k+�އ��o.�=���@�%���I�6���}f����#l
i��h��vd�x!��F����"���wOA�s�"��Hb4�"�'S�*v�Qp�L7<�9�D��@|�gF�
K�p�'�.����R�U}�?$'�n#J/�S�J V��A�N�H���n׮XbB��)�8|K�s��D�=C@�v���F�Y�{�\b�Pcyu)k�M�kB��uqZD�E�k����D���5�֣62�<�U�-�~@&��/d}�#e`��#Q�L=~pЅM�H�.e �����egr���@d����F���4,i3�Z�w ��J3�9� $}7�;�NБ��������x�~�v%��5{c�ϔP�/3�����Q"	'�-ĈqVΫ�e��@?�%�;7�� �\9#�?��9�S��U;�a� ,�)]� h�l�[ �՝� �( ]w�H\-*�vj�k����	�����0pņ�+	�j�ZU���.�1S�w�%t���!*���J!�û��2ϲ�Lp	�aD�T�!T�n�����Բ�N���H������te�f='�*tL��f����)�^��i8;[��^L�ŋ�'*����ǅ���}?�C,�Tw�1��M@�jMr��Tf.K��ېJ��̀��1�
{���`p��P��jh���ɠQ�{���[��g���Ԛ�Lc�>7K3db!��ٞ�
�_<Zw�����$T̫�_bj������ՙ�؈��cGLj^��-�G�rzWcQ~0[78^���}g(����#%Z�����,����5"ĄQ��SO��� ��R�,�A|�.R�����(�"�՟����,�,F�.�7@O
��㸄8�I?�쾩a�d�{坄
ڞ-�!�%�Rވ�9?(��Q�;Q��~L���]�\�#��DM���{4��AY�V�x���2%B�آB:3Ҭ�;���N�� �1�Ȁ��@�WL�^��a�JVO}�����1GȨ�6��)p����`E�h�ś��F���Z�����ws�Gl�h#j�y�n���ʯz�Ό��3,ԛ[�0�#_Ƕ�j�5�%vkq���n�[g� ��ó>��������M+�ݵ�����3.��?��wE��Jɂ?�R.hZ�t�Aޢ<y��IG;1� ��=��Y��Z�ui_tpc$��t���o�����G�њ��$/�ΞY�1��"^ǒ����;�~��#U{�(0�?�7��`�K�vUK���	+���ű6�;B�J��2|X��
��2��k�5TQ��䑭*/�+�GCA�1�KÉjMVSM�bH������4�u�K��f�ơ�;�=sGeI6�*5�R�`}����yQ���I�x��+���t��L-H�`8���I�bi�b����l6�O���A5Z(�QSE��0���K�6��&�9��A�!��gINWv��xn��S�M%��z�>�ݘ*?�ݤ��]r�ݱu����cy���84����֜GbW��d�|���sĐV̒�*�_"S�m;��p��>î:Z��Jr�	���I�I2�klt����Uk?��'aÐ�#9��{�89�[�k����w���`s�9�"�>���p�5��J��<k���'%q�r�f��8�V�@�"�Q����b��Bv���w�:1�8ڿj�)��=���$/��b��'ᠳ�����݂�U$%�f�H9]3'jx� ��R�=�4�}}�Ѵv;79Y�$���ƴ0���+�t��g��e.k��b�5�*N+�������h��;h%{��]�EO�BD|�(�T��O�>6�f���on	�^\��SN\zU.`����E��\�dy��� �
������v/�[��51uRxl"�˔�o��t.��+��G���j��(���f$&�,�X4n>D�_�x��N��+3*x �ْ��s~\����e�"��ݨ���0o`���m��+oH��фYyAV�����?��U&{��5:OPj�+̏��>U|��x�3�ivjZ^����!���?�5]{})��GE�[�(����1@Xw����q$kQp1ĽB����!��̐ZY�-d+�7���2ݑ8����.��Fw�V�N�Z���R�Τ�C�%"�4l7#��# �7����C�����c�vي�����ɞk΢� rWE�9+"g�ዉE5ս���z��Eg_��dm���,��Ĵ!�^�� ��hM9�O��}������#�rG��̽�o�C�H�uyuHV�*+�g2�8��}OL2���.�=j8en�=�6Bm����Џ����c��)5�Χ������䝡�FUm���b�k[��:�;��|6��:�r�5��#���8�F����\�(�<ٍ̀�#��>Ǹ������J�Ʌ3��@�N���ϳF.Г�{�J�=�=���&��wL	J�vAT��&IB�-ĥk�d�������h�&����1����g+���,�ڀ����ƨڙ�U�KO�����]�n�-�皈g��7"�4 1$3�ޅm^�^�ŔtH-+�,����\J�RS����_T�&������U��}����9ǂ8�x����eM+���v�4<���d�`в�B"�M��p�SQxIҥQa|�n<�%K�������N`<����'B���q(���"j��2&���<�9E��^�	~r!Sz�˾f[�}�b��0���Gᬖ�|q�Qf�fT}���%��@�xW��ҜO��x���hҙ���N��wY��d	��}�%�ei#nx�hP;�[M�ۇ���Vz[^R*b"�U�9�BȮJD�ܜh�6ʶY�~��2X.�_�tW��E\������5=T��V6�6��i8'�����D��1�(n�dp�}��fak�f��R�����:ڇ!d���zCni�:�<S�Y"�'���*�����
�G�~��%F$�\5��LJ���0c���f�n)��\nT���}q4�|��:�g�J���pû�5ݤ��.!N�ψ�Ti�&6"���cTN�TſdT�1	�]Y���P�m���;�|H�����Zl�&�X����`|�iA0�� s�9�@�$-�<ceV2Z���q_3-�� �'o�����;��}�xp��|w[���e�=D�ݲh��濫>�rƤ��F%d\{��}�/�6�TJ�ф�$A.IV92h���oU�ݥ	���Ф�Q��"�P>����Bn�2�ڥ^t�������@��������+�:�a��"U^h��Q=[�:�	:B��gEq
ֺ�X�S���iJ��Ƈ��O��@N+!�j���oT3W�{�@kb���	Xl�����X3���8Z�cNV�Uw�Ό'�������r��eӮ���s���ʃ~5ͪ*H���j�	n�~U[A2��'����ez XA��h�m�Țg�ߌ�_�9���I8[c�?�sI,�nɟ�	�Z߬'y�4�����$�^7G�A�ѩ}�k�Ƶ�x��e�>����d/j�����\�4���Zٗ�J��}7f'��O� �����^�`�?̺g5���<�(J�v-�����G!�_�I��.BR����|�[i��%,�e�|�n�+jV�8�@�X�~�1�f/���>}�d��k0��.�~�p�{!�k�$��ږ��xQ/���l4 �CǕN�u���ug�<SH�;�␿�`�bм��moc���
���}���g�|��7���RJs�Nl��?bL�M�~�ŕ�m̲n���S��1���s���aS�����R:�o�&~#�G%gʦ}0^�%V��:Z��Q��r��1��?�	Q9�& ����K9����FSaR�S�72!	���W�!�qaRQe��n���Zm�	.c�*Fcb��=~$�]��<OKV��j�<�T���׆�t���OR��vȀ���7�#�ʾj�&�W J<>�H�J�`�b'��#�L�� ߳	�w�әb�@mKio�OT�����<֥A��V���coE7���o����L.����z��ᔭf��������dۊX�k��7z�Y[��H�\&v q�(ւ�����ݧEK?��TD�Y�Z⊅���UeH{&�U>Y�g z���ث� 4׳VU�Qc��n,UVF�e�p#�z�93�~�s��Κ��}�E<�b��v�4ݿ��^�<	?R�S�1����H���Q�@�s���/w!�~���,����+�b�8���'^^�� �<],�B�%%�w��s�"Y��b�$�⋢v�a���)frK�-%ۊ����Ul��PRۿl�!���]�RڊB�3�������
W�X8M�K8�5;6︚Y��b'YK���E"<�7ی�?�X$.�U��
�u�,jtdy]���tX9��sE���z��XiDA�X�G�
��g���S�fa�ͪ�n31��`I%ijU�;-�/���/$�n=+v�&�p���C��\*�r^@^0��B�D9əM����c�K��;O�-x������;��V�3��j@�5�|�tU����M
�E�"C��ޮ����R�����'�H�\Q�r��զLu�GGPT�$�WD�������{6HB��o��y�R]]u@���*݀~�)X�9Pk�<�K.�g�@� Ή�P�b+^�ncF{ Ʒ�/bj8���_�Җ�l�.���MP�$�P&5x����O�ѓ�-A��S?��_96:�����6ߊ�N�LK�t��CK�W���I�N�����o�a�t:ڡ�/�bZD��@;�
r!�jk�y���7��N(X�9q�c~��B ?�2mK�ciFA.D�d�/K�Th�����B~Y�&��(ݺ�8��`�O)�*S����H�橼{� ���Z�B~|�yŉ1��o9]�'
��72���>�Y>T;4@�%fוf	��#�N��(�c騗tC!�4���F�xN~�B|n~ƁG�ݐW��E:=�P�ة��)7�ޚc�x[���,�`��x�Nq�e�6ˎ�h���I_����x�o�@z\��6G�'&�i����u}�q���*�\x�����/�ף��*��s�	J5`��vQY�Z�)z�:��涑�]�F`�j�۟H��.f�]ڶ���L�!�e�c3¤Sj>�J ��/�d�X��o�V j����#a����2�����ςk���Q��a_��%�gp	Eh��葆J�)��5��&�\F�gX#V�Z��ܣ8�L`D/�Y���H�w��M$�fv��&/�7��>�3�1K�Sɉ��b�
�D�1=c�E";�+������M�$�D�� �q!������ �p�?��l��nE�A�]��č#���^�>��~x�ɮ8w��,Uh?+o_٫�X�j.Pt��uc��"����Al���3<SRo��2��^����B���E)��Cu�a-
{Ə[�<+j�(�_w(t�7���t���iē��4��� �����B�<0�����hx���0x�)R�rG����t����X��Kx�$��U� �{1����9���RF�Eu�{"%�Fn��C�@�4-��2|\<��"`�%HKwQcq1�r�;�m��Y���.��7 ���3�󱛕j�$��w|L�0�W}�����D�2t-l��e~��Vt�gg�Vd�i���&=�z��3��yId/F��x#[r��x��F��c������JQu�X��ە5>c}$��#�p$_ʜ;J�*�`k-v�=���ݘ '
q!q/���ٜ��5]��RFY�29c�9����J���mq	K��dQ<Oʵ�&�39�cn���:�iY��`1A�ׅM��ݠK�m������pq>���2������P�!d�-�$���_WN�h�UN�CD�y�H4���h���:g����{H��d1o���5���k9��z�Z�S��e��{���}b��k$��D"�����dh���=P��|�@�[`�k=��c�:�K�����GfI[��4����#��D`C7aTo�F8�\��E�������&$&Z������h9&��>'G