XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����O�h3$b"�خt�ŭkE#C<�FUc�d4�[�
'�Q&��a#�(��T	�����&쯘<��}[p�Or�#�p35��O?`��b7�;8}�*É�:cM�>��36�)V�A�Ϡ�� ��B2�����p���-?Bbgp�,�S���3@È��E�߸%�
(T�Sf�k��H�F�������ؠ0ǭ|��Saڊ�N,��0���=��=��)l� ���rt�R��vA�ӁOb0�&#�Z?�� �[���Z �b*����q��o�k�Jw,�V�w�n�8z>g�*��Ӻ�	H	�J�)�&c0�H�wC����bg<��e{t/���
$����_��r�##1�u��.\��gz*#E2���:zU��e�`�X��M$��&�uV�y����\��mA�r0�uF&(�c�u)#�J�K+��4Ș��!�J�cN��ZE	8�%�>����^=/z�h �m9)�1g�����4ҡ9;�tw�Âh������l3[�p�#�}��q֤J!I�7Nf��\1Z����p�$��;�jr(Z�|ě#�k�P/~�0�>6�HA�h���6�!j|ߦ&!�^���h����O���ɴC+�UB ��'
���Z�8��s �E��p�M�3��f��ѩUF֊��8�$���Y7�_��!�q��� .�:5eF���ЭfG��(7S������*�xDPt��˸H��E.�L�f��ӽ����Xj�R⇰I:`�+�b���d��	� �XlxVHYEB    1661     760D.c��)�1��wi�O��-�����_3%����H���67�n3�[���6�)}���f��"���-�����I�֑��s�hu�����-�/H0͓SQ@�<γ�Ѭ*�k˵��ֲd����HF���pX�9�ל�>����E�Џk��r�~0�i��7�bti�,���@j�*�L)���d�*Q�^$��S��#d7�q�'D���;1U�Q�'�8�7xtX�c�3����}�s1����{�!%�]v�sH���R�LD8Q���U�H��^.03���ͥ�EB����TOw1ߑ�(�y@��^@��)���7d�eV�t!�r�s� ���PTT`g�Zk�EgD��F����
b������� �0�u�H`��>'�a7E�o΋a����5�;m�d��4�@�W<k��:�բy+K{c�r�f5��;|������5�4x-Ac|w�y��eh����v�M}R�R�0��e>i�޽7a!�&.,����M虳���jC��$�V�>���S�o�N���Mc�u�3���T�p*I�r�(mE��m0	)e°&<��7�&U��ع3ilsi����������e�Ue��t�<7��M��E#&�[͠���������,n�R��B��eZ,CaT�"��VՂ�t���}(�Ա�X��ݵ��Ϻ�@�iB����&�5��5d�%bΦr=��4OEtt�b���C�l��lkħ� 4����5����!ѺJ��j�b	C0#��ƼLCG;Ck�8"�G���v����OΈM�{�ht��ؑp�>{�
tA�c}�/�,��L
�6p�b<��=�Be��?v�Ӌ*ؘ��x$4c�q��ʺ��1�$#���:�,Pj�:-TC`�o��#~de�1�T沗�]!0�K��dTαȷC|jD�� ����ɻ<�?�:��%�m��~��W��Ȥ�ķN�����`�����7�l�1�\��o�&M3�J11���s)Pcn[�4f~�ۘz���v���We%�meӑAc�����N9/�Unt+:>��x��Mb��opw� v�����_�j�[��~%��}5��Rk�'ѩJ@���W~dtU�����Ybҕ�-#�M6E�?*s$�H/K�O����R�<4����4��ܔ�@����G�w-/�Ox�*&T ��#�h�����M6,ur�� �`���o2sL�/k��[�� ,(����E�nB1�K"@*�	�|A�����!��Hʓ������X�0.-	��(�e�I�e�I�s7�\6���oA�A���x4A?�n���*X|u�ڭq��b/��[AE6�Ye����3H06�Y�����2�G����R ��KgD簀�'��Hx
v�U3�-sk��v�Rֶ�=nы"W_a?$$o��V_�<4�и#	����� ���ELX�s���hVQp���6k��ҿ�a*߷��Y���Tj�? *Ϡp�q�@�5�� m#�#|S&wC�V����H4��Q�3j=�a��Yd�WgH�=�֣ꊵ��yU��1�n�������i���s�3�ZI1󩹅流݋������5 �����q}C�Ĩ8�(rqp��L$o���栐�vK��4gvݭ������ُ�7E7�6c��E9A��N2��;�2�޵�ZA��H:�HO����	�wzp�FC��ʦξ��+$�G�,��9��g�IВ�`�������ξ9&���<���B.�TH*�W�1-��x���*���j��N�Uj`D�/(�
M����мSi%\�6�(��dB�w2\������H����R�[(�>*��lc�S�=�z�\v�\WM劎�VF({����S�2g!�����쿲)�u��