XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����o��B����v�����U�Y
�]���'�'�z��v�޲Ĥ	�&IC唑��@��*�y��`>����]~V���졔��[��M�����O�yqC�}ص7V�����R��	�g�<
I̵�s��NҺT��I��<��L�5S2Fy���d`��9����+oZ���չǹt^�X�B�W�)�r��c�O���2�V�r6lJޘ!��WjwսV;wf �^�PH��l���,��YO,���t�i�f3�v��h�'���ja�$g��G$ߧE��5�7'if4�w{������k��ï^�5�8Ң��:&=`���-���s.)~�?��:�vG�]⇬��t�_���OAC1�� A��$����<3k�������	Er�0)72!��gw3Y<��Z}�
mA��oF��<7t\K�� �����P#���!�rb�����z;|6�����)��� _��y|�
�����$1?J����h���.��g���&l��C��26HJg�)C5��b�T�X�K٭�@��L���$R#�����s%Z�Y�m�����<�BK=H�z�=����?4����H��!�� 2<�ŧ�9�PA�2]ӑ~|��+�ɫ�E�~Fo�^ v�)�0Q��������a#.5D�(;H�;I.���2�B�#�F����R�͏2�C������Iy_(,2s�b%	��@,��u�nѶb�p���S�kA�z"FҨFXXlxVHYEB    1001     6c0�'۩9����� ��C��'�L��|j��)�}�d`w���x��w�Yq������� Ø>�i���>Ml����V��;�%yi�n����P�8�1ű��Y"��wl��I.�P%�|G��'�{4k�7}�����
W
���ɘ���Qo*�,:�8�O%Ļ�5FY�Wb�]�����5�@,i���D��~C�	lӍi�p��钹6ء��Br�-��I�΍�d��6��HZ�{d-#�i��;�/;s�c���ܓ���%�`�`3^�x�h���Uu���GH$��P�Q�=
J���/�V��ɆŁ8�f�����7�ܰ;�W}3-��d�5�qA��(XV{*��lCۂ�^lT7F���Tb��u���8���C���x�-�)��,����i@�sN�����Ɨ��r���w���-+W�����NK6U��`�1R�;�jT�V(�Ys�^�O�z����񶡛�$_:��%X$���y���+hIu�v���R�B�O4E�&d�~�4J�"�%��㖅ߧ���Z�Y�Gc"���#��(�����J3��7V}��Yy��%��Ʊ:����*���ʜ��=���;j+������&��D�������b�Cۦ�of��c��x����׻Q�E]Z}�z0�%B�����
 Ƚ.R'���aG�ǚ�=�����OveC�� ��>~�`���e���y=��}��7��)l��O��ng]���+R�?��}ӿ��	��b��,b�9A{a�&�o��_7��B��.�n&R�/��k����B���xq%���-�YkJ���͔*��J )����r�+�%�	����Qe0���gR2'��}���0�F���v�
<{
���ت��}����Jc#�0�b�:�ԏěSn�>p��˚+�r[ :ظT	���̑���WA�-��{�vos��C)�mJ��.SO�L����IJ�q��ݭE��B�`<�(}S���ڻi�Yu�-~Ӆ�P��w�u�sy&ay#F����6'f�!�P��:u}?g��$/��%o���ѫd�.������ 0`2��r��	6`�AMg�1b�X��.�"�˨��NrX0��n90��vcS���lS��#����.׭�jK����<�Z3ȅ��;{�zO�ݡ%RO\r]�@P(6�= S���5��kZ7x�<Z�:�m��?v��w��l���-]�#�{���Fh�4���r,L�Հw��a�ֱ�l�0�������1A�g~��Ԁ��dҿT��\�Q��Ȏ�����am,j���vՑR-7�P�p ��ʘ�YQ�"Cm-��="�Dv"�@���3���� �7�1���f�6��SN6-��_O�y-fd-NHs���@A�
9M��vRE����b�V,��<�k�7�c�e�j�-G]�$�:�5��YN)��+y ]|��RTE�zѫ��ch�W�����	^�4���{��>	S^�MN�Dյ�.TeAӶ����_�N��j�O��m�-}7���Å�Y��s��yJ��Qh����'���51OE�RR�k?����e��)̩�8�ʜs/�&��4�Z�������u=�\> �M�jk�r�T��;^�[��Қ#)�>��vbn�3j ��WJ�%���7�P��2V�(����!�����"&J��O��)I�Ys�~,�W칒G%�ߕ�_M�­�adB��