XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����]M��|���#���{+S�ҝj���/��,4�y�Y|���..Wܑ�ZHߐ��;���� ��ZH֗צ�,�דff�ׯ�/�8�9�r/1	ӣ��3�N|ô�nY�W����6�$ S>�
�졊6��ȵ��ʓ��ٙ��+�"-��V��ٷ�����a��'%�U�j�m�ϛ��W���(,�I8�K>��c�m\���gx��~V��w�$���e�2RG ��s� O�����GM���mR��W���S��t%�\���J��]��*;����7��?X^���F�^��_�Q�a���&�g%'��!�:X3dz���u0+�a�?��Jf� ߇�ة�|l�R��<�R�C�5�Hk<e��E������@��ǀ��3��m?�v�?~z���:#�A/�b0��'�V���a�| -�I���#q�Ս��]o��Ȑ���ȁ͓�l���Ue�ے��GC�`i��_�����eq�ʩ�'�V��.�ÉDH4S5����o��Ps9�τ~��&���X��G�4s�cNb.��#`P���42�]_�eظ����I�����.��ʢ%��0Na�W��k\���w D��y)�'��(H?�i����॓��#�3i�2�KH|L��4U&��7ia
�@!����k�Ӱ�&V[�?	� eV^�)@�b��Z!SH�j��ݽ25尮���ޢ?{7K��)h/��j�ŝ��\����[�ҜF��Q�W-�(�s��z�`�g��ߣ_XlxVHYEB    4071     db0�YŬU�[��4��c讉t���i(��� S:f��K�ݾE2����GY�mD�.��Ԡ��ȼ�I���:˴G�6�!K��0�0fnǒf��������r`49�]��.t����"���$'��mЅ؎���|��䉿:)�	�5�dچ)p�ǛtN�?�c����vj�Q�bd
�U�9�*�2S��%ߊ普�f|i�v��L�,���,xN�챼��m9���[�2���.7�&����L�Ҥ�⟊� �L��H���d�a���ULц�t@�xF�D����:H =Z�d�7��,���M��̽�-�m˓׶By֫����wq�f�i#�;)�VL5$z���
�� .t*�(M2��E�Z��f�4ܤ�`��5����1��>!7��Teg��t�����;��w<S���\�=i�,/�����1밶St�NX?.'����Vۄ��q���%�a�c�!�F2ܠ�����!������m�n�5�_-N`�D�6<����?7����U,i��ub7`N�4D˫�_�Z�(�ҵ�@5U��ju��D �q�듁��Tj� �&�`u��r���Z�j��"�k��גag�����곶#g���!�h�A�G��k�}�K����2R �Č�|m\��nɊ�|����ꆉ��ez�묡4c���n;3ɚ�AU�G�C�E"�c����R��&��.�Lh7�q'�l`�j��]�C��ۜ��>�e�ɲ�Ͻ:����{k��IB�{�O���ɬ~!�\϶Z�3���K\
$3��L�-�| ��&&�_�RS��k%F�߰�6�8H��~$_��X���,��;<	"�G���y���v��g��M�@ވ�-f~�5T��\�ZyS"E=/5�*�{2���i5������h�����0CԙT��ϗ�p�������`O��d��Ї�%�Uܣ7�PB��WQH&q�����m}���o��7���^L_�<�E2)؇(k��!x���h�w��F#�b�M�Ԅ�˔��fnI�Z������Ȟ͕�q���ے�ú�>�e|R�"_�t�h<�bקկ/�����������_�Ѡ�c�x�|ρ���L�+Bo�,����K�.�	`4L�"~H^oħ[�t3e{�+�xń��s!R��T���l���r����R���3y�U��A���<�s��<WT\'��d�ȹy���m;�A��)������$�<w6��3[�9�w⟉�a�_Y��s�������m�{���6{6��`*K B��:����bst���rq�<X`����25�ጐp}? nhh�=<�&���$R37�=�M22�	�Q�˭����T甠�P�yS�j�^�,Yͩ����.)�Avr��$�$۟`Mth|]�_V�Y��D��!'��~�QXr�"���q끎o��Er�������Ȼc��AHC-2`{�.��_D⩖( �K�ukK��s�"�����z�R6�ވ�&�:y�����j��y���t�7����k����A���~���3� �kï���W�#����VSJŔ��d��Q2������9w��k��8�vZ� �����	��}�ǀ֚��섊fӚ��|�B����&j>o���"뺇¡[��W�4-�� j�#��(X���Q�cd��C(�P��S�g_���(�PĔ�}6������VYo��SZv4��Y���]W��E =�� 
\ͭ�>�&FtX���[rxwˤ+�k�s���@Wp���3	/��tc��R�OM�������2Q�Ja�4�|�^.�όH�\F��G�8oТ�H���+zwd�$���	�-�<\T��5��w��S���s�&Ix��(s�n'��ްi4�������|�������*��v����Xn��V�p����Rx*m�[��b�'��*�x#�g�;Y$��U��z#
��#���ԡNHF���B�Qy�a��%D��K5���v�� Zp!v�+)�XOr�,H��l�ҕ��";�L�3I0�$���������������5�H_y��ܚH��;H�wa���h�_�(O�Q�|���p		�r6��"Գ�j�[�4c�I+�  ���1�|.�˒�R@���F?�ft��o����;�[o���M���M"�7�i"���K!bx��E9�S�;�uiCN|#��N	����k�k ���AsO��rE�w��+�dכ�#�չ�����aU�
�����Qwy�k*�q�ɤ��=Gc'ӱr �;8n8�V��*�2�zB!�w�ý�>����xRg�{����z+i��F��ܔ�k�E�b4��n�[��j<�$�/�^;�
�B�R�^COlo�� �[�9'g�yn;��z�(�sΠm��90�5��8�"���Z�\�e2-0�
I�"Ƀ{Vt����Z��Hܣ
r�!r7����~ݒgp6�u�$2�� ��%�ӿ[�垇4yh�䟻���%�NLp�9�R��(S�4s�e�,����:��Od�s�p��QP�I,��2��r;�
�
�	o |�$�`�к�V��I��#�w,ҿ"��&�{�C����ˋ�o:���*S�0�[�N�H'���n�ч��n�9��$3���%t�٫��A��,�X�v����N���׉ ����A}��G
'��8��lh#f��lX�����w �82�YW^�E�8+D�ҧ�f�Y��%�����uB~}��8e�6�H�K�^�&�C�Ι1\e��a��uw�t�D<����e�j�
E~�e�ur���8{�ج�p�6�X��tX��nB��d��p#m�_��߈P��bd�R��$����)���0�#q���/M�Y}n��I���o��ڜ�p�Oc*'���-�w��ʖ
1OԜ,��a?�ܻ��(�����|�F�B�_�b�{6����~���O���|�f�cV��S8�֍g��%s�#@��� U���[�7�.D%&��K�X�ϧ���sg���+I*�cȘ�vM�+m�dB��/Q�7������z��`m�X&6;,Q]+.�����ǉ�m��>���g]�J���/�Th�N����A�b�$�Z��CH��:�tG1��.O'�	B�I��y؝%f�Hŏ�*�v�<f�{�r���K�(���-z�����I��ӝ���2������p��;����WZi[��E��Lr��F�q��tǑ;�j�P����~f[\I� �ʱ:�O������B^X ��|�wܾcFr�֞�=��w]�vE���(�,�l����s��^�ܰBT�OC�,�y@�{����\��'��qQ�,c����m�؇�;&rTO<���]�ߕ" ��qz���6�q�r��5q���91W�?�zg�To0�Fh�^�����y�P�HDW��|�c5x����	V���=B��eL2'���/J����I	zo�D