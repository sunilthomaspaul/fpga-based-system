XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�� [���Bn����8���}��T,��`QՆ������!��&������[0c��5�����7�!�"ջe ������]*���i�T��n&8ѫ'Oy�|£�������	���Bƚ`��nEH|}���&���,O"~�ؽ��̍�}l�Eܩ�)&3*,��B��!�����j������n�����@Z�Ŋ*K�<u��X�"Nۣ��`�l&���-Md���%�~��-�hX�.�?���n�wJ:l��>7�OZ/�Ҁ�7iN�"h>F�i���EJ�&p�� ����o�sA����p5��9�5mg����D8�����e�����_ۦ��G�CX����LS�h ����ƍ���YZ���<2��NyE�͋��ݕ华W�{�~� �/mq�X��
?�u�E��>)��0�$�����S1���]����7�bn��:i���-�г~(\Dו =}��Z��X��'TǗ?:H��.�8�ɘ54^G��!����¸9�uuo��n%�Lu��c��͊�2��9�@#����I&ߘ'��]�<Y��63<�1H8z�}�{N�>5��.���H����
X��.���D�F�ܠ��5�[1U�{i����WgAhI�h
��6:�k��t�-2S����9\� [�Iŗ�p�~Tɔ���/8H&q��pby�\R��N�|���&�W�Q,]�#f�7��<�D&_�."�BK�!S�Z1[��"?�;�2��M�
��[*���"/�?�s�rXlxVHYEB    3f19     db0[�l�g,6r,��6�rʡ���6�H���JCM�a쨼d[���vO^�
;�/Sv`�,{\�u?�f\�}z��^!л"�N�=#�M"O}:��ʰ͟���܆�V+Tª�BF
��s���w���#��Q���Cr���x�20?j�e������懹HG�n{��H D��	`�P�א�Q3t�gq6���#I�1�i����Ǣ�]�$ P��
K��{J�1\^�D��1�0�I��7ŭGpB��6���e�N/_���A��Krc���B��b2��ZӐC�X�M-���/�� q`0���h���t�P��D/I�-i.�Pǫ�r��e�� ؔg��������1n���JY6���rK��|��nW���͘��t,�t�9^,}	M��<�N�X2�oܾ�����f�q�|�����DL���0��9���:�L��a޽j6��䉗ǯ�3�p�H�Op��)c6�����F��4��I4;����r�������g�&%Ʃ�-�������vQ/&	C��Rj,�����;ΣE5�)�Dp��K�`��<|��*{���^��e�9���	�.,�j��4IXuW�:�t��=�c*�C��rN�+���	�\�͑*3�1s"!�rG8�!FɋEE
?������y=�Z9���ҵA�]���!�-������	{��Ur ��l�OƸ,�l�w���uD�O��P�*��!�9�����������]W��Y�u��|�{�h�I
cU�g?���6����%]����4�s@?�qauf�p��=������Fj�@��N~=��G�g��C5����q�?l~+yJ;�+����[ԍ�^᡽S�Е��ܤ���$�qi��&��X{�&�����qЀ̷���fF�Z��ƫ�;�	?(�-/�8�>��P�DЧ�-�D�� F��2(����bQI	�ʪ�t�G,:ȍ~�k+�C���.�i�Xq�Ho�c1�|�v�wS��+��_^q+��ʓY���1�~�w�>X�F�mj��o���$�����N������ )-7������XZH:�LA0���|�����k�%�~��*?��C�`��o*������4.��Bhpi:��,!�Q�$0i{e55r�]��T� ��f��D�*C��C@�ȌB���U/�Y��7MQg�W~%ye��[A��ż\ �H��wT��\	�6��]|I%]������h�=s��@����P%����A0Fæ�{�e�`J�z��lq��h�v��5Q�L�s�B�0-G�fdx�����!)��U-�Z�����Q�R�"O��y�M�}2�BrBE��h�寢�cT��E8s�Ҹ�j����c�;n����1	��ѝ˭�V�f|%���jR+���"���'V���x|:J	A��pO-C�Pfa܎ة�p�1�
�t��.�<f�:�o(��֌�O��8�*쇯P��Э�ϑ?�8���^n�/I�d��O��4��z��I ey�
$m�>1�w���}�gK�J.>܁�@�{�N矹����c��(��d;1SHm�d�����7���A�#����ŭ�68��.�%��
۲F�3�XG���=DߜB�u	�T9s�CV��ѠdX�O%q �~Ȓz��U�z�t�J;����;彨�e���~�,դG�B@�;�E���	�u�Ђ&
:{�i�|�.���"�ݔ�`�v�!����u�р�$������r�޽�}�7I�)��+i���C"ŗ�w�H�[��טp�0�-}���_C�
��>]���8�?$>*�nb��IV7:t�&O�f .��]І����G8�A���8�l�5HS�8(dGMVj��V� ��;���1�\�r���ԭ�~��T��F��  ����^�Gӱ����_��).}T�]��P��� ��9)�ո���(Q�^�$��hຯX'Sj��#�#������^SY&��P�׿%��JcZ���,W7y��c\0+��w���A[@�Ȩ5ga�v(�E������	|�aL(]��avT74�Ŧ}꽻�&C���0��Ҿ�sk��	�x괚i���+�Gieذ{j5s��Zf��+����'�r�L��튑Ւ)\*���"�h]�B=22x�ӐS�=&�B�%�H �^O�����`Վ#rV��B���D�y-���f�5�KA[�-9\�I�yO�#�����*���cL���-�آ��w[���o�Q��=�����;yƓp��D����O�h�o>��Q�"+��f!>S�F1�	6���8Ju,
�*�̧*u,�"�yS���N�^?�o�@���$�6�oz44}qQnZ"�]����\F�� Fr�i%�?��`��������wn`1d��9�>М�
���@�A�#9�>�T@~|?Yi2�c�`;�F3�Z1�k'f�������Y���t��|H�T�QKc�nL#����v���g9�x�������Ǎ"Stc� N)�߈FIG���,������M��J�:T巠��^��성�o�,P��o��jg�|'�WW���3�Mu����������a-[·en4,|,&���J5�+6&7t�CƖF<��Ԝ�"ہ�Z�2P��E%ߑ��59E�Dn��F��;a}���ݱtC����ikC!ʱ\�܀��;�r�!�c�~=`��ɋsS�V�k�/=�|��P*�m"���E�} ���G�p���<��n�eU�<������1bĒ���#��xM��2}8SW�vs+eX����΀�����ajJb�$�Kc~^*,�YM�7WA�����U�Q�2y�L��~�{/���x(���Hh�T�ϫaclM���M�t���.`5�p�� ��U��Z:�Pz�* �O,\�\��a���xs��#�A7̵���Y�hy�$)��[���U����= E��&���_���#L'	��U�5lct��ȕ��K��o	>���ؚ. ����������f4���-\�loE�z�>���V����Z�ώ#&[�a�\��/��ڡ�@W�^)ݞ��,��տ�mh�7j�^�惾>����A����e�:��r�p��T�]�?�^��W���Gf��2�n�b�d���U���y�l���m.���d)��ֱ&�ްc\$����H�Üj��s���V �<�H<�n��ŭZ��"�Cyi?Fq�4���v����\D�"��=��~�}e|}�JY+p奙İz[����È>#!�)@v;�ؗ�e(Нf���"��@�8��7�O>����9��� ��[t����g��-�
�q�n�}_��;�Y%be��D����~L�hphI��y�(�i���b]P� c��x4 ��H"��WH��0,ſC�D�|��XzE"�%	�SՁF�����'�9rLk��~������W����v��1�2o+X��.�Vӟ�L�D��(�!; 