XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��T�G���wi��O(I��҈T�1PU�C�'�+��r��O����1K���`�Q�nro��;פ��_+��2#�CvO�y� ����_a���V������G���|wbܡ����N�k5��4�Rm��B�3�7|���p���9�&)�A��/����\�W��,�ਨ���"z��̝z�0�]���,��",
+>D�w�z����鶋Шd�Җӽ���G	殉�78{�.`�v�8�.-�їF��"c���sL�A�˩#��h1J����.�d=��v�~T��8����|Ua+����!�7��d��TD��YA�Ww���G�J����>r�-Y�� ���H��|`���ig����j[x���zÆ6,�Pl�%٠�*~RwUP� �l�����Nl�Ɋ�L}�]U��4��D���%"k3��擀�_�TK`�.ĮEu��J �����{���_.h���UT��ȱL�&{�j����;E�Q}�4�EȖ��?�tl���;]����~��6��K�&)������O�DZ��ƾ��������Wc-�?G ��l��,u��	B��R*��|4��%۵�L�84��{��]��)�D8[u�#:��@��Mꥼz]�no=�w�ҡ��X^Y�Ƴ��n�S�v�6��Ӂ)^}�3j�6P�G,[(z��6��2���y�{J�(��W�%�J�m������^\��y��z���83�:eJ	���bjFX�XlxVHYEB    5fd1    1710�v:��$V7]��E E������X‗yAf��n|��*~z�E.��ބ�t����ŕ���#�7��R���5,]K�p�����n�r3�����D�ib��0&;�DQ���H��9��w�W��^�����j3��f(�5�%�E%�x$W��L��΁f@�,�_�ꢠ�7�IlwS i���g�u�n!*j��o3f�ME����N�I�d���v�M�a�%�;�B+Ex ��#�fB�"�]�4���a�����{o�)��6���/߷$ɦD��V��!8�4o��ѿ%i�r�����M��[�e����آ�J@5k�R�|�_#/Vr��|��C�#��<
؞��kU�T3�n^�]i�Z>�y��|"��^�!��$B�n��ITIدώS�`��W/�+cw���i���uFrhc��ʩ{��M�<����0 ��W1Ӣ���20�7��&X�\í�䂫�O�e���X�+y*3��c�Ӆ�MV��9�0sRɱ'����n�x�� �u��
{��i)ei`��q������/�n�}�Fz�h�����y���_��	�p��u}-6��s��r
zZ�l��	K6����*%��u/%�F���p������~���+�|��U�>;�|�q.�</� �M�D��R*B�(��{�t`��$��9��3�-�Un�V;�-O/]�]h9ut8���&	/e1V�^��=�*ᇾ9� ��
'�F7�p}r�\���i�9/A�	���n�#�����ȣӖ�����\۬����Ca���ɀ�+�F��'�ֳ�ۛe��fl����Gl%z�
�q[�����܇� ϰ�$\@)��q>��
�K g�R@��LA@���*���wG���M,QRR|\-�h�����u��a��I9v�#6F��O���/$d�ou�?L�J�N6�L���X����yv �"ɖ�&�]'�6���ߩ�I����#����c�mH�x@�)�p)����ɂ�x���.����3q�+?:'fC�-_G<�/�{�I/�n�{Ĕ ��)�����h�mR��X��d�J(�>���eF�Q���9�g��t�A��ώ(y,x���������y�/WG��3s`�}� ���)<b!�օ����a?�E:>�+<{d�=wW���C%�O�Z3���;lAv�Ta�T��،5����^�eub!�G����|#�B�{�YsN{�9�����{K���w���~�^���F%0��zT�U�
W+���?�@�)�4����#�ҏ������	���j�9�݋��
��Ӗ�tp�ر�[}��"k�-bOo�1E�]����#���J��^����W?F�⪒��t���������\� v���x���a���<|_��� !\�kצ�L��i��`uQ�2J�:��w~?�N�?T��L*j]לj�^�����&� N�˖�C�N��t*g�vR�07m6�����;R�Q{�p2���}�Ƕ\�mx�������:߬����떇�D�����a�c~h<)���'��̆7�4���$A��\a�:~[�����Ffy��e�����*0Ŕ�-��`H_����R�*WlӊuR�?j
�V�$�$�RŜd&�ZgTJ��ْ���QҹB�.ir��Y�����m��T�*+���]�R<���"e�ǧ� Y��"�Uϰ��Po*�*6�� s�	��}�d���������\f[��c�Ǔ5��W�*��PO�q6�Ȼ��G����*��n��`9�`HH���U����v>��L�
������p������Y�)�ɨhW�d��増�=%�ɦ}�|�K�{� <��XA��$
�j����E��h�e��U�!��ΧcM��T�ez�Da+{�~�^��><
vm�Z�j��'�zϭ$r�|
�Cb ��Ր5)��:Bv�lV����^����qV�p��T>�ܞ��8�kQ��P`�\LKh���Ep��`U�!% ����Z֤��G���[.�T1�-9�|4�	#t��&TP�iMX����4�Qpی��670X�ˀ��D��v�'�-mY�g�C�	^H=[���y&PZ 1���F�%�R�bA����m�r��\Jvy=[x������v�0�u�G�>�/x�
�Ԏ��5ؕ�t�w怈�·����o>��q�vO�Q`ى
������޵fX�Y)��5�|�7(���{n��z���p8G����Gڤ�Z�2ݱӗ��0��+Tzm,���0�[o�dJ[c`�w���J�P	+1�3y�5��HJ˒	��3��쒸��2�}��+�+e/꒗�W�
&��j�� �]q ���F7&d��.(O�f��Y.�:�ɄP��B�o�Hه/"$Mn��V������X�;�ʯ��ڭ��6yt��c�޴W�SH$�tg2�H���R@��[h�aⱊ��C�)���<�����4���$'ڥ���N��	V��@��h�vζ��1����Q������̃�懮p�̸H��ޡI��'Z�;wn��},�0���?e ���e��	�(UtB�<��F}u �,��_���up��e��&Y��@3'Њ��_wI(� z�VV��J�3,QM������OB(�Ъw���SDsqF��X��~��naV�.\+WF!���R7�z�| m�Q�ˡB��F�a���!0�yC75���I����e�4����C�u�ͣ<�$5r��n����U�<q���d���)�ݑ�Y��9;*_�����M�Ł@f��;�.�C�)�������C�n�P�fKϥ�xm��Y�zG&�pGOr葉�(������%��w9���\QÍ��;f����~�!s')yF���R��_�2���L�,_i���w�At�����.E��_q��	��"�+o��R�R_��@�uV�7�gVcVk�@����ӺY���/� ϻ���(������OsZ��f�_��s�.[��$9: uᶪa�a��O_׋���ߦ�S�LyxMi����˾��>���y�tܝ?�]YM�d�ZR���k��~ԯ���n�Y��������t�>kƪM��6����<�8� ��s�15EC�f8����2����5P�{+,�%��ͦ�Ňۍ��П������jW�Z+؉����wAÈn8@8�g�No��{`+����A@:ZPE K�3
f�r�>���ُ�d�ڜ⧛�s�j�	hk5/�!W�1>�>f�º��J%�\ǩ�B=�S���#�
�5���FX�?���[`���m�h$��R	+����,�r��ް=-������ �8=Ĥ���&�q
Tof�X{N�-����5]�P�Ү�^϶����A�Z�KIuW�T���T��A<le�BýW�M��7 �X.[�/���&:�6X�s�)`�E]�G8���H�K-}���B����<�P�\C��4Ƀ���X�9q����O�9ǎ�;�^Lk֚`���n�>Zy�{v
P�r|^��
�����>׸H	��_��}l�SJ���{�n��幌�h���a[N���E-��%a�y�}�	��W���YM1�I����K��D��/QT�qng�yP2�D7��)�����%�L�M״W��Ã|�����/�tK�0a���_*����!6R����E�Ͱ�;���ƫ���� ��C�;DV�IB.�6[����%�k�+nW��98�LY%�9�͛���nQ�r��X)�Dٲ\���u��WJ6�џ�!�%
�7�S�
몒��\Ơ�Q��f+��47�9��෠m�{"b���!9���"ʿH����T�'@�A�7gM9w��'p�*�	4O�T�L���~���^g�q�H�h[&n�o���A]��G�!����s$����?�AYޞ򂽇^�0�z��fw���`�O�[�^���g/�2�}�S�m@�,���0�i��G(?����/c�9� Y��w��p*�`�������W��hw�)�>� ߈�j���H���4�uҔ^��G6[�u����,��Xܞ��()D_�~Ŋ���؆BR���FW�*���}$Y���>�]K��%�� ��^���pL�5'��JjAtúݶ��B�u
0�������I~@`l�o�v�5A�r��:��h\���<�Y�d:�dW�ӥ��J���jx߭NR���3߂2$����e/�K��k&�P�cZ$��o��Qj����#�n���(�M��7�x ����[܋@�\�D��'�/�Q��NA�Z ������v!h�|��<�ݴt͐IP��NyXHsx7N��]�QOR���5�$|e�w'�I��J�
(�̴��<[{�$��w�9N����ꮏ�U�U��\�,���" r�����%bc�x�.a�Uw�=�+�A!k)lM�ȥ�U��k|�]�\��&���@�c��o!��z�[��V�����昀<�`,D�į�,����8]��J�K���l�Gp��s;��s�5��L�h�T�1�-Ƙ�����W�&x����Փ1Z�+���C��U<�ӭ�@ݍS��'�}�p���Qu�Rg۽l/:����À�ߩD<E=���J�5�oL,���]�ӑZ���f��p~M��G������eU�Y���ƥ
��w��83)��1�ՂiO�V���?��5���B���^��}k���%v�>�Y*�Ę<8��x�cB�OVK�R����M|�̨suK�k�����y�� f��_D$_�����n��B�F�D~��å�S��]͓}kA�b���Dts1��<�Q�hYo��0�Y�l>��DS8k�w)j�̤ loAh���� �W:g�]���-Z���M�;���!T�:Aiz�D�;vB�۴1���'��'M�`��8�N�J��1@赡<O`�_eXre}�]�Z�ay�e�&@	^?pu�\_{���!����I���e�!'\Pen�Ҡ��>*��aDc��a)�Pj�?��9FP�N}��R^��墰:�x6�/���Y��|_�3�*���J4�����6�i��"�,�B�u��*y`�:�tEb�.�oFQ�Q�ޱǝ]�فG�gt|�4���h빑JG�q�G�+HJ�!�Y�\e�����\�$A�<Ȝ%�'�(���kv9jꤋ|A�7���Zm�D}Q��Aj�t��L�2���l@����e���y�5�;����dw�>�\���ʟ�R�v�(<�K���*�k�֍�NQ�ͽ4�8�1a�u���� ="���V��T�8q��'���BC�l�Ρ�.}gm��{8���" �b8�������D�V�i	B~�4�)�|��d��U���f����t-f��=]��fX�~봉��Z�P�jJ\,4�wי�7��L��$������3�<����M�6�������wF�I��P�1Z!�[Y?�E5�ӵp\q�̷��s�i�uu�@~$?��i0�;�Ub�e��eȄ���yz},�RY����Z	� w.���-(���Խ0*���h<�@cT�:�̚�Np��G(92����6\$�AX��w��� ����k�ϖ}?P�	/;Lˣ	'ؑ�sh;ұ��.�i'�,�v��s{���.bv�uk�bydy��/����4F�8�j�J󈋵ڷ�\t�!�+́?�rZ���\c�{���K�F�#D��Q;%�IK��|��������N+ɿ\����K��U����|BuG�W�
0<��H{4���'V�:�!��)f�$��B_D6�j�R