XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����=����n�VBW�`\sGyH�T>���~$v9-��	%~8t�&�L�xUe�q���v��#��t��dM)��蜘���;.�%u��ރ�GG��r��Ceǜ"0w�'�,[Y��{�@p.%<�N���c=h����x:݉}	^��n �baԘg��m���	!��|�$��)� �N��ݗ7�y9��1d(��vw�f��`�H��lz�ao������> F��β�,���!�E����D��҈��!���t����	O�	f9ȌG�d��o/��f��/��hT;S���H챌�N�ఔ8�,W5XV<��p%̭FWZ��q���ն��2r�t�̀�w���	B�U%oX�C�$[����վ����w�Y�����%ǯ��`߀�Lw��R3Y!t��K(�,NS�^@O��'#d��P���?���$&1mH�����ƶ���L)V�J#��A��y'�R�)���	���	�m፵�c�1�F�B�lX���9�03O�d5B�Sޯe��41��:Љq(C]��$-��dG];st�+^�V�T��j�G��q0���\�5�u�eGE �J�B�Ԋ{��T:Ҧ�Qo�z������|i�?m����6���HvU$V�p�(k��N�*G|������_�w��Wڢ�<��� )<ᡄM2&�B_/���˟иUW��l+_1|��E-�?��S�#d3���Y�'����&xj�O����
��lw͂9F���AV�1f��9��9`���ΰ�sZXlxVHYEB    47d6    1030A������КE�r�sf���Z�$������D݄6�	�kg�WB9��������ht�	�Z�a>p���S�N7Y�=A(vL��*��d&�n"LF�h�0�nCۈ�[ͥp�w8Ó'L1RJn�+�@�s��9�샓`}�K�v�������"�L��^�N
DT<�$W0����V$p�$��V��Ϋ�t%�'҈?ſ*�K�:��?�[�$m� �sVw��+�t�/�j�,�x�i� w��~�� ���>�e��^�f>�v���R�(nY*��\z�P3l�N��3�3W$��"-G�~RKWљ����&ClC��^�Kw�&L�.v^�ݻ�� C&	�D	��<����<;�C�u	!&H;�w�
�^P&�.1k$r�Ԩl��?&�a�Y]��HcȲ:I����la�rݦM�e3loK��io�ҚX��Zbr����m/lzVn�<�N��7
�?)�����`�x(S�N�*R`�?o�F�{���9�t0_�|�R;.A*TX�kXzk���Dd�~�u�J�/�$r�v���wK*-��-
_�  �>U|y�~VqHof��.�C�����N<ț��G�7C�=��+��M�'�d:b#��B~��G��%�ʮ{D��͇��G�4K�@?�����%�"%��;�M�V�.>��»s�i��W��q��s5ɔ�@��y���g��1��cs8o��m�k���zz�u�&t�J >��D�ªr�V�m�$�׆1�&{��&�����F�k�%��K1�ik�æ���16L�*�w�q�V��i���DIΑj{r�R��\v�B���N�����E�c}[�e���EKMX �G8�5�sod��Lbw���TC��T�\��v��l�!<KDj�z�͞���6+ې���v��a����[�?a���EW>$��:C��|Z��h�*��^��:yw���r��T+|0�u�!^k�J�~�%�rC/��"�S���/�g�="��7����׽  M\b�o/
�x��G�l2�?�\洔�<\�ED������ɕc=�`�D\�'�>Fy{��v��0+y���d��I̹txu�`k�(`J׏�v�(�B'�(4� �<�^Q�P�����Y7z��e�|w���#8�p'{ӏ�f�A����L_(�O?~����!^�K��i��Q�]� ![����^��J��3w��*T*�(xO�]���N�v�����d�:�D~�W�\�:®t�4�õyx\K�Q��� e�m���䇊P�Z�v��mx�W�+�F�ZA����(g��q9�
c�&v�1"5���mD�����@E����od0�3����Z �S�"�u@`'�Af��L�_�o�m�w���#W�RLɬS�Ps$H0oKC,)$��~o���Gn��Fy�͵��5��p[�����G�㣣F������,�=��;�rD��V%eyi��n��7��%�[8�C��-n�-7Fn@s�84�A���P2���lwrȃzv�8���B��AtDSS�x1�����EV���F� J�aE�"�uc���:�X ��iޢE��(";E
wRǝ)A�0���.�L>��7��R.�K�~�M�Q��]ӎܧ�n���%4��ȶ�__�Oju� #������sUb_\IZ`zVu�Z�4�d��1O�|B���sӷ�����D���i��%��h�>m���QE�y�o�����{��aX�������į�h��2�&�J2�z�K�P�&��
W(���Du��t�ybe��ћaJ��_�?�#|8w�z�/.V��[���Kd�<�~���
�)�Q'|�!G΁\W��sT�w����b(G �a�w�R!{��e
�,��W����'�|�F�2j`��CP¿�s)h�K�N�7������U@#<��fd����;�N)��>_cӱ%��0f�v�_�i�q�/�EZ�����S����9��	(F�c����h��^��-�HK�u��M�ŞX겐^�^\�h1�YjVΤ�eC�l��-�����Qiq��TH�/�#}E.E�+����_�n�����_���{HpPG�}uj������R_z6��S��5MP��(���G,h����י��q������iv�`�����1Y�
ur��=��:��|#�X��5�3Kv��H3O$V��	ک�ōogC��5"��܊z��㛙Z�vg�g����lIMԽ�<�bI����2���"Y����P���@�P���d���g��5��_�J�JF�p�%�|r�$N��!�5%5��Ж3�\���ד�*�?�@#&�܄Y���#�L�RI�.�&3_S��*qA�H��(���p��
a�	�c �T�����⩝��S#:�r� �O�A�"H�����F�6">q������2̫�BMŎq�{��_����ɤ��q�p*=9����^.��ʬŠ�qT3LHg�n4���Dd�1��4�@���<|��N]�+�}�O��%ȱR�j��AkQ�� �DI�"[&����7��t�9�_��f�&|�>�7�:�֑�9�2_&U��I��L�c!�(���S�Q���%z0�H,����}�>�v�&«-|��Q����̓'MV�Mq���u����`6���:��Ԕ5
�4j�h�V����W��P9 ���?�5�k�N���@/�=�$�䎇�<3�mGV)	L���a�k]-�̇t�P�c�k��|���Ym�!"p������1��o��#��e%�����'c�˃c�#'�H2�"r�ι�A�X�s9/�D�471{&�O�w�ϒI��S���]DWJ]�������E���z�C�Φ����5�m(WCDh�;]3�R�bJ�U >��Z;{S�5k�vYka�ú�u�.B�����#uS �Fust&ٰ�х��q u���7����ni�|��E[�!�OQ�0¿��G�o����K׽��&m��.����p�g�n<���q���;��I���o���������v�Z�r�����+j�L���w��>�z��jlc݅�Q�����J��G����_��;�S�*|1��%;�W*���K����P��ڵ�Gz�ޙ,��/^F�J�z}PnjEJ�K��X��N�蕜q[���Zn�j�{����Hƪ6r�3�ہ�o��""��Z6��%���\V����u�GC�Nw��[��*x�Ƅ=�P.���sO8&�2�J�.�.}jE�|ib�vB'��^/�E�|�xcC�{�~7B,�Q�u�sbEb�_e���X��?Oe�zipO18�5��?e��{y�e�G�F��$�L�b��B�ӸX�Vz��t��O����YGF��R�e��� ����~����"jb`kz� _5�@��,sJ��U�.1ж���K�3��e�/t"��([<)y���s
a�ƞ���I5�����t���mMk�'�N?����E{�~�p�WYe�!�)tL~��2?�oa��bWi�}�s����ݪ��V� 	��q{{� �%�Ědpu�5�Vi&Ո�	H_u��.�^Y}�W�j��VHhq�f{�-��vC��i���ea�oq���.m�V�aT}<�1;(6O��<q�BPʹ��C
�ߕ�Zz�՞���
m0,��Qf�
�˗��T!�~�`�m������;�!�kO��d����1���dV�ֳ�^��b���0�C��3f�V��1����r|�=�����ջ��UpU�V�q�8-�*�)v��&����Nn"���VeV$Зj�8�cɖ�B�4v�o#��f��m��hu0�I@:?�2���%@T>�M;�l�*;+���|��31��<�+��}�":���A�O���3�v�n�`5tp f�G@�`���Т\�4��d>ױ�d/�ir��M����:0I{1��%�Md��+R���;'��Swz!�)��ag�(�8�r{ܲ(��:�<8Y��`��ۦ��K�`��)K��N�������\ȧr�����ۻ����'5־�ތ�`Ta��$(���Ͼ��ɌRv�uP����w�^ކqEc[�IA�0\�:jN݄���@��*�݉X�b