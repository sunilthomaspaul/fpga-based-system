XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���Ł/�K��L�,R�{��|ٻ;��@���	/�*Lul>�4��0�UcǱr���5m�˛��zG��񆟖�K���|�4.����?$2�Z�:�c�C�P�j�SQ�N���;�x���fK`#�~#Sj����s*FlsJ��LV��t(���y�Q<L�{)�rA�fj�8�5k-����w��y#�e�,m�2�N�ti�:W���L�K��qk8�B�^�Hmu�x�k���4:��~�`^n�#*#DNP31��,>�0g�v"l���kL��� #w�A\@�?-��|�^L��y��s<^gM�x?T�����2 W7����3�7ԡ��>�|+_,�O�@'�@��i�q�0�b*W��I1l���Լ2vY��2�Gh����~� �޼��ٜ��-�p�g�ʍ��Deߤ��hg]6��g%����_"
sK�eS��޻U�����YEWz=��ؠW4BK;ǉ��=��o�����^�����p�I�����F�5��Z�S]����J��W)m��G���M��? �+8�ka�����g��NG��������y�zFݗ�щ�A�I��R��O�����azc���lZ(\'��.M=j[��:P3?x&��Ae��ƯՐa}T�v5tN���o��R?���`�l|��2h4M�-���l[��yOF7H�
����&(M��R�h�8�v���ib� ��nY-4�9`zWpM+����"W�\r�q�-�E��^r��XlxVHYEB    159e     7e0}����dPj�~�R2~<�4�+�G�*i���m���hn<t���ݩ+�9�6\���п� ,!�ǡa<z�Ώ3nv+DSyå w#���z����Z��	�o*g��O�1+WR�%&��jם$���s��1�|��Qh�e5�!!5�}Zk���|x<����,��Fw�W�����؞�38A�Z�f���;@���&P����b��t���go�C5�g"R�p ��&9%d�P)
�&�Q���n8Zh#�N���њ_z|�<��5'R+��F֍sH�uK ����U<w/�G났��e����p1���h�������9:��e����"��H���f5���Ď������{t���m)X�~�M8_u�l��_��A�U�A�#��4�w���l�f�s�FtfJ��dr&�i�9��>�c'1|�&���� ��{���'D�������j�Z��o�A5���j�z>�L�@T��ɰ_Wt=�\��7�'k~��4��2��/�}N"��G��:�R/΂�	=fD�'rp�6^h @!�1)������
;vQ�y���0�L�Q��Iuw�� �0���w�M��\�-��;�����a����0���k&0sjO�d�9p����)�����
�.��aZx"��t58T��Ϭ��fh�:�C�v_x�AV~}w^� *��� )J2��n5��WX��c�\1�6�-{�k���b���5���k�۔0[�.�����1P(�+zj�6HfL)X�*���Y��,�Sڞ�����w�a索�=��Q��������.Α��o�<V
�v�Z`���af�P��;ʿ�D��y����)�k_��^�ɯI��_��w����
A�Fh�^��"��\{E�y�i���Ui���ʫF���}.����P��݉j.������Y��VD�
1�,$A7���ӛ������\PV�7���1�Fz�Tūd�=V��VԂ�UGhXt����r���iyղ_����@�A�L�V}	 ��/�=�K�p���i��eJ<Ѐ)�	�?;x(���V�)m���<G�&u�y���L���*�ߍs��F{�2uu+a�"��;Z��:��-���?<�YGi�~Y�}���[���p��oժ J\b��L�9��;�|���,��f� �	���ϋzz�ڜ���▬��~�4���"��ZK�:\�D3iXc�8���ɘ�����ې��*�R��)H@�i������ͣ���[��:biN:$> >�m\�&�%��p���3P�6�Z�������r�a@y5�S�}��OԖ<�àWQ�l�d�$q��������tL�!��@d�����2MK��� Z�~�	��WH���fR�|2�Og�@bnAa�fV��E��v��ф̶%���3���M�x-��z59ҵy󣟼+dW$��f�=%X��z���N<-$&��y�M��z�>���,�Ֆ+K����pb�4~�U�m��K���q����^��}���pB�:�f}�^~�5C�=WT�C��OhZ���B���f3<�J�� �d�w\�Q���l1\$T�,]�B��V��Y(yݴhׂf���2c���d$S��\��,�Z�o�F9��`�+�]�2Y���v�7�^\Ogې*�9�HM�Ȱ�V��|6U�K��h]�a�[
�5����3����܏���a�u�&(���IU��n ����0GU�M( Yk�7�@P�X��f�|F�Z�a�?:��4+{L�VK��,�� ����䢒(���C��}/�I~�E�D��g;˚h���s��2r<V�;_��$��c��#A�R��'�q��/�	�œî<"ެ/�F�����vp~5n�}�����L��iɑ�l����%k��J- �H2!�^�݇{4r8HЦD{�1��r}����nU8K�r�0�9U��P�%wʹ��	ٲ����>�9sFG��v��Q�����v��A��������