XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��ؼ�O!�u0 ����C�a���)��v�������7�B�y�\���nm-�.%.�I��F�1wZ�z��t�/̈k�=����|�
��cǞi�[�B��Fǅ��m�W_3~���ZF�a��0s�"��K�"��P�b4ol3ΐC�fm�� d�mO+���sd����6�7s�2oL���k	d_|�[_�Ez��	ØX'�s��	�~⋜<΋�~�#2|��B72��_M�7�Y������-�j��q;ؘW`c��A?["xx���]
�1���n�ڵ�g^-.�җ�L�הּf|L*�TӲwKy�����c-�1���dﱕ��]ՇQ9h-�aKě�U~��}L��r'F��߿cU��V�μ�����V���w� H0��7y��9�9�j[Q�ט���-�P�G�z�SS���� ��K�/G`��I�>�xl��,��ݒ�I_�$Fu���_���O�I�� QUm�`Ѧ� W�o�����i$h�v
��������z�u_8��~�{W����	/�C��Dl�b*و�ܕWB�7����x�B��~T���u��_0_�o���	ٮ�yk���#+�?fn�p��!zk�?��EL��>���u�~�߿h�s+��B*�: KX�$i}��e�e���yy�G��ɲG��l�s߱3�5h>�qX@ �%�Yh�A���!�3Ӣ����H�4,hT���g����YAo�MZKg!Y��ERպ�gG����v�^�G�����U_���XlxVHYEB    1001     6c0#=Am�vsJ:;�c��5<�l;�[��m�!9Gt�/@����EyuUP���g����g��.��(���m�R[x}����+D�娃Po�q�LXs�+���u�	��{N ��v��Ԕ`i�e5�$�0��	��"���+Z}���c*Stk�㕬e��sZ��������WJ�i<��7cI���c!��u޻�7�����9���2x/��L���PG@M"u�v��-�S�KR_�PEȋ���c�R�����]�cmN���ơh'� �@F�?�����#_F��{��}~�8����Xf��:(RM��Ň����h0��x�0[�Y�ҳ�]��Z�d7���h%�E����Xm��fV�)�4��V���S�-_��:��I/�ך��e G��D�S!;zZ�wI"1!��AJS�.�=W�*M���8�&�^�q�D��;�tN���A���&a��8wH]�,@�JB��U~Ё��U��|�cP����&��8VXl��ٽ�6�=�&D2)I�j�$:�fȽ�r��q�b{w�f�uo"�����B) zB�N'�=��[�q�r��H��b�7�t��mA���������IL�Α������6�/	�R�3D��L���gK{��D3|�HDl%��@4�&gm6�޷�j��`��	�勰R��tI!��w�5CU	����{�Ed��rx���[��i*So�}�6�
vaM ���S�s<�HЖ� �^��5N�7rۏ�*S�MW>���)s�:�����Y;N=)S3����,�3��\M��_1~�;��<�d����XA��3�8�����T��C��1Nf�aH�r�d=(C�O�F@�&!�ˑz�{u�3|lI��A`Ծ�I�n"z~qةU���	3�k�u�${��JG����%�L��8�˶�7��c*������ܾd�%�n�
�,_
�A�s3��O�ќ(MH��F@OI�L�����ۗ꼘C���0.u�:0��׫����w��9���H���8S^��MI�s�p���[[Sk�!E���,w�ĴS�̛C�t3n��ī$�����g%Y�Q�)����ఱ<`^�;܊8�G�ȝ���;G���u���2q4r/��ʹU���ƨ��j��%njv|�dꛄ�,��J�O���O��o!�D��V`�����@C����|�R���W�d8�[͌�T2!=�m�O��,%CK�[�׽� G�Գ��´� �i5��$����I>F�M3r�0��lS,q�-�0��c�kb2M�6*�V����ڀ�b�<��S��W�<'̊�����3��1�2r�}O���G��':AB'Y��^�B���������_�����=Q[$�QƲ]I@NO�v���]qYZ>�q��+�'h��\�j)F���`��U��Iم�lr���^�+\���L���ʵ$U���#0�D7�'^����j@,���Q�����
���9�p�4�������[��83�+��� �Ҝ=��
ʨ�\9k�L�.�,�[����걼l�[:͹
R�A��F�9O�7�]�"�O1�j�p�1����C���lC�Wio�8ݤ��WRy����WЫ�m��Z\�z��N��V/���6�E��F��|��*��~��e��'~O$ë��������4��-OL6P�5�Ģ��ZOl�U����<H��ݼ