XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��y/-K��p�~�d"*��e���^��=�u�_'�T���{����U6�AzssB�k��xf��*'�*nn[S����-�j���v�����Ā�X��[1m�Փ��?�/�3��
��b%���L�������(���7ZNۏkx�Tj&���V8�4�0��i�� ��w�0��1��,߸\��҂��$�Ċ�l^zE�f��C��݀";�|�kci��wzu$���f�/���9L��"�d��mqØ��+̺��2�F��5alUg�!o�|F��7�1�}�U���Tsym����wJA|���h=9S�km�$"\�W��>j�GVo��K#�_��5����U4��-pQ󓺅zc�����C|�/�-4�ʽ�(1�R���� �L�� �U Z�]�N���vZ�-���5n��9�z���0�NYe��o��W7�{��<���yye�]eK�죍N�s��0.�hԦeP�n#;W��M��r�k�>��x��ݓ�9;:��t���a���5�E5v}�?,*�/#t�K�5Dg�W��VM
ԥƾ�L�4գ��ʽɒ�9\���c���e ��tz������7�"�S��+���&�q/P�@�)�\��I����t�ణr���^���%�2$�����WL.�����˧�M��:�"& Y��m��~��b��,��8h���)�.���~Dj�|� ռ�]\��@�P�d��[�I-��2K�|�i≈�,`�$|�i��_�ӊ��5�XlxVHYEB    1231     7c0�׋��J���/�+�㎁b��O�.��u��?Ti�6h��kB��Y�@c�(�(o,�4S����ꂖ[��)���)�M�y�nVg%q.A 
���y`j� �t�;����Z���8]��zl՜z��5$�$���Sl�����EQ!�U+[4-��謬�ƫ�Z}p��rA,�C"���"��1g�)�k,4�/��0i߳��R��fmL����,#~���lB?)b���y)���CH�%���a�>Q���¿Zu��f>�$�-��?�$XY�+HN�!�̋�j�����i�>�y׶2�t�%X���#��RФ4�8�9�Π)́��63��3Mp�Q_2�{;P����Y�s����Op&����B�C�3������'('{�O&9����$S��+O��t��K��Y�o�D6|�?�����й�5����pm�B�-ڶ�%T�U����^��o�n~
y�;�P$�L�Ce>C���,�h���(�D�9��O4|�؞�������n/�ib�����]U��r��J$����%�"�0U�v��E"���Hy� \�%T?-R�0o_�5�:�,��:��H<��lqק =��G}�1��{Ȼf�W��T�܏��բ���V6�%>~Os�
�߀4�c`�Q�'��4����;ҟm�3��=������R���!� �e	.��#��� ���'=�|�T�h��b3��E {�WS3���Ζ��y��RM���|"ۼ6�GܖѾM�V�_'7��*���#�9Ƴ	su��J�sS�soʮ� �=L.*=w/�9����g�In���F�i��4����@M�� ��y���Uȃd�/� ����ϮS�(մ���4T��|]<��i�˸� �&B23r�q+�I�<��7�VEWlAt���S�M��='H����R��ݚh�{� =��F��&�Pȝ��i�*83�Dj��~1��2�����Wu������ۇ���iޤu��A����_>7�r���$��	�ީ��,�Nq��X��*c��&T=%G p�.�'��?Zi��"�:9�2��-��j6�뀳l��Xi�"�)7߹h2D�^��<Ҵ�jԽ��� 	��[	�pè�Q�NP�M���ˊ,�`��>�ɕ܎�����|{���Ǵ:�l��f(�	4�ty%V�IFgi�ŤP�Խ)p9oR�j����ݖ������D3��zM��	ϓ���*�9���,�L�� ����;��:�����KM��l6ق����Fk��i�5n�_�l��o����p�� {�d���N�_<E�82a
(��
{�A��3�o��`��\�F��V��cQn�����PB��2���D��_���_)I����P�v�o��`��1.ŋ�}�j�q�E��ȫA�s�b�3��&{D�{�P��ja�9>�&����D�J���Q���a���:���n�Lf�I��L��X�c��.����h���kP��1֓��	mT��})kY�S�wܬ�L���ڈ5T5�\3��Ӫ;܆T��"�*����?�r)�7B����p�������aޱZ����@�lD	%9�x���p����A�%W��:7�w�n(691�
A�x�NגN����Z��1:�36Lxd
]��M1��0���ަ�J�� (6<����/±f��^�u��?;tYF`:#F�"f� L�U�9J��~��q�О���ؿZ"��(��Bݲ�������W�t����e��;���A ��6jw��ʶ���.�Eh�'���� �n�EbJ��(�T��oN��
g�� ���Q����H��� �Zf�X��//f�ڡ��;,�I���/�D��|؝y���*�����&��:�B6��jv�z#�m�8�Sɡ��)�0i���?�����{��!��Js:1��zQ��>�6��|�% ҄������R��WQ8^,���