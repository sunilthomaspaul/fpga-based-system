XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����JV	�Bb.�m��r�G)����o1�<Dh�i��*��C��s(�yeD\]��%��s��0K+?V!�������87Zb�|ӊ���'͚Q����9�j�q�:�ET)S�ٍ7f� z)����i^����q�6��ɋ�c���H$X��^
��Px�ç�4M��"���H;��q�e��G!��\�á�7���Dy�w���+[����&E]�=����,�UVLf�����WW�Ѵ����y>F�ʊ]�G� 5� ���搳�IL�![u٬�b�s�œ����x�Z#�f|�{$����Гn�Q�j7�P��+�~գ)]l+�r���n��iFȎ�5��:ɑ7���H�>����~'=V��S�P�Ǖ�J�b	W�@t3S����і/�S\� C����"��q��5�P�j��NPTh�YEzCr���5d�+�G��n�R�T2~�A��jt��Bpӹ�}��[&��Q�ճ7B]p���@N����@.���e�<�L7.�nt�ăY]Y±����GK3��'N��<�\#CO>e���-HS��+ߔ�p�u<�S�>0�����My���ILՠ��Q���#�Д��h� b	���P�)�wG>�X�ݺ�
^l���)��Q��v�ȁ�ԁ����F5%��e�!d�<��?
��yH��
^�n���9�M<���>��.U�G���d�Sp9倎���������`!HuO�%�Pb�%cOM9�*i����tXlxVHYEB    2fbd     d20���'���$=��m�h�u�k�/�ˤ!�'��݅��	����ep �;�].��D,p�p��Q�lꅞ��LS�
��CZ�j{S��ō��M��	�@��.�~��<G��X�����C�"�b����H���`eBT����Y=�*�&�����Fxep���ǥ/��젛���Csؕ�g�ߊ��Gy{�|��kq�j���c�{�/�Ƹ�˭�]�8ڶx�%"@�!>!}���07]Ʀd߂�h��?8Nl+�)5�� v� �]3��1WRY�S�/8i�`�J�#�mZ�U	�Ⱦ'?;��>҅�zE�Ú��+������3�qQ��6��.��q���-����,�@��\�=l�/}u�&2�[������r[��l8��pĬ�5~� ���j��Gå�\�o� q����L����I�*�.j� +�/����Pb�&2&���4���l�:<�l���m�X��Y~!�B`tH��'F �����#�_�_p�q/I�r8B)���tA�1@�ߠ�c]��kyU��tU����8�^�����h����|$���u|��e�H�om�c�˼ZB*Րӄ�� ��&�f�Pub�Y�2b`lJ��6Ԑ��,|��TfE)D���ҟc6,n������������
y��z�� 6a*�����b��TM�z�dv�����k�60��>�H
f��w�v��Ȯ2�|�Xn@�Ȕ�8�n�����W�v�D�9��SY�bT�N�!��΍�A�$�_���,9خ�k�N�����4�,7ޗ��w3�
��)-�
.��!@I�j��H�ld�TB\v�_�����<�X�|���c�C��^~��`o�F�3���2��&M���OSHu��4�$��$�y"
�B��@���ï�yI%�ޒ�h6&|���1ur�N�0��E(����"���No��©�+�gM��	��{w�ba�ַj�ij������� ���ѧi�/ao���7�����C��IMF4�I)�+�ʦ��˸�LW&u9C��j��[|��w�����~���E��h��$v�5�W	��"r��S8�Α9�f�����̹U�ISl���B�+#�65s�?h� �n#HbB�.����m�	5�;�Ŋg3�5TL5��c5�%=굮Ӗm�[�x�h�Bs����3B�m����ɓ�h�4��X��������{6�t�?�&�=��]�*ior1�-�����&�Y�hL�^*?0��9�"7�M���Cd��<Y9gnU��qy\q����Ɏ����f;�zڡ��M�.4J�ݘ�v���ʚ,���VÏБ����%OU�>Z�î��4�4�[�P/�p+�Q�襋�-Ƒ]oz"Ɂ�~�49�zU�I��椛�?W���]�{�<��އ�o�dr�3�]�r���/����I��
��[�y���R,Q謑2��mVî�d�1f��K�}�m��t]���l��k�5Sg�ΊRhlf��g�E��OJ ��3Y�:e�M�������n�P�k�Bwr�ȴ��t8\V=��ϖ�c�`�P4GO2���E[��w曅�)Tm���n�q���]:�B��J����\���S�`����Z��yx/�%ĴU���6;�m�MF �U�)��-��wǏs� c"�� v]3��X����;*i��!N(�uns��4�C�$����ÊrOvi�����
���C	6�X!z�{I�i[���1�hfmK�ߛ�c��U�������(.BY�>�S���Q�k:R8�K�c�ӞX��6��ʫ��݀����8w[�m��=��t�g���wB�T�b4/5����XR�������VLH_ow�[0�+�>�߂Q��ۤ?GV|���G77Q��/���$	�O���Z�$��;%�*龁]��\Z�ǼEȸ��*�-�����R��"���.@��OY]���=�N�4�]Uh�·���+"��X���q�y�	[��`�( �L��s|`4�2@��I�
"��^���t¦
��*�ޑE�2䮘ʓ�^�. � �`�U�T, y��U�[ <
����V�+�E/��P�Ep�=jF�(�!�J��x)��k��E)@�eە9��M�?�{�u6�F� 0IƓ�@�j�+�b�Tah���G7�%@����e�8����I����W�д�Q��	:��&��b6&!�g��DDۂ�U��T��ឺ@��If���f&����Q}��W�X�?mRU&��� ���x�P�q(�,M���V]�U�;�Xh�q�K��wC��F+�A}�mK����yXK�aU2S��0Q~����h�]J8]yiL
�<�E�8c�aG$�F%7yJ�A$y�!�T��Ü ��k�Q#���B֪s�����bw��,�c��}аK�e�CZ/�KQ!� �O�\O�~Ň�z]��M�q H�������E���K'3�UM Ud���ll1C�#�=��,5H2�[a��?���XKeϛ�oUC���C�6?���$6���:��	�ל�
�����z�}�D[$<1�ey8��l~ @�{�>�wX���a&/�i���p��o4�~ ̇������E2�z�	ƹ6yPy�goG��.�f��q'z��b�ߥH�����p���c�Hy�S��h3����Q�)�='=��(���ڬ��Q�>�_��d$��D=�߁E@�)���y�v]����{	����.��@��`[�[W$�Z�!0U�ڂ���D������Jo�EeU뿽��&��0<
0ϣVz���'*t��d(��^�	�`�*MYx���	�+;;]�.�O�?~en�Œ������Vp�޳��3c��S�I>W�G$�V����Z��Y�~k-�3�}ڻ�v��?8y���_�l`q�ƸY��ͤ."�����h[��"�[�E�}Kּ*�8N�W�ѸUXYV��6a�k����Ƹ��fw��P�Cݜ��>r���W�c|��g��0,6���P����{��qK����
f�L��%������VG��ngt�6T���<����4�(_���[�ײB�Q�=���q$)�>j���{�r՚�*��'t�<9X�0~��p��db�l�IHA�=z�ՕNoA#|A����k�?�}zc?@Q�rpE���:0W�ύ}t���ruA��J�F��}6ΤHyBPhӳ]%5�_ʅ\f��\������7Z=����wYnQ�yE*ir(��=v݉O���?y 8�����o�e��%Xs�h<�