XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��� /�2vy+=f*+?�{aX��K^�X��y�L@+ԇ�V�Yn
m({M����}�f���`���v��g.�"?�p<qT	���T!�� ���uWX���G�y�u��ఈ<3o�7�#{T��o��ПY4И[���|����j��'0���B����̞����l�F�# ��t�$�׋�Bp�D�u[�׫�Gs0�3�Z"9�X�K���5�Q,�	t��ι'_��+���㪛
��͆��
.��/��$v�*Gl?������Q)0as�����I�`���[��wq%��h�c6?�H��Y���W��0$���r/�E�v��1/�ҟ'�9�_j}���.��H��\kȠ��o_�Q!]�A�;/ C��ic�\yGn�J�E�ˀn.GhѨ=�[�(��wcc=�|Y��䘕|�2��K���r@n3�=}�uV��h�*y�t>��\&�IL�@��C���|N灯�q���sY��o�R�E��:\vK?�m[��
n�[ Ж�^��e�ۀ�N�B�l(�6X�,�)e7�KN�x�-O��f<%���d]+�M���mZ��
?�;L�{V+�6��{#9̼�V�|{_8fMw��F0������=p�r ��
;\m��#�bj��E�g�=%�/_�p���t�+7��`2���L1�C2 >FY���<Y1�u���2��Р�شP�±��)@>9-��ʲ���V;��qK� ��n�>��/���bkmN[���M�M����~���XlxVHYEB    1d59     8c0�V$�� �e���HA���f./�����fC�cN��ɻ3��5�8��0M�k5Fd�,�T; �[M1�g��ڔ @���.ά��I/��4�X�`I}�P�֨f#�@G�_-Jo�L�/�,˳�eA��e"!�.�HA�G���4�Va��m'Rs��n4��T��3���Đ�\�թį���4�ӘG���b���}4Yd��|��[.x������"S��V�
}�LZ`�I�x���D�}�h�m�}��=^J�td]���N�R�w�h���Bw�XULh�*��cEi�&Zꠤr��NS��3� "8�y6PB��<ؚ������)퉗[%{Rp5������S��Y� '2��{�o >n�*_�X{�P�b������%iO4$eΔ��+�{1�%f��ұ��k�%�׎U%Y�#���bW�c��jK?1�����ǟ(�S�'/�O�mI��2cE<_OW�)qs�i�3�>��Sê��$� ���xR_#���]\�M��,���`d	
����t���������+u#3��O�953���%�
d�*�%�-�b
8�6��?�]`�Iw�:Š��Ǔ1j��g���Ϙ�X��&�H�����m���J�B�ën�Y
���-N���]u���ĺ���`�򵔂�z��.�h��Q^��I�o2�#@��m
a2�}��b�\��N�w�ɪ�1rN�eR��i�=��l���s�g��T�p�K01�9��|�)B�q̀��o��r�#|L냚z�7��R��� ����P���<�J�*)ٛza�{ƈ��z'�9�V-n���O&�_�Ɵm8e��,L������`=+���dw�����Tw:��Ut��l�_�!��H�_S���g�[�=OI{���� F�$1yЅC
�5	�Y�� 3}i�
�
X^��Y��<p=���Ba��k��._	�`a�Im�� �V�JL$e�% �y��{�X7��~�"�
�P�g�TC�U�����z �';����:�Ǘ1����i	�騂U"�.ɹAO�fѧE���?%�f�DAױP������򄱬RE/G/߰:��J�}@|O�.�uq�`+EI��Ӛ$n�H :b!�[��R�Q���2טi�ͱ�_z#�&��s�a����=����n(3��c.(�+츎l"ki��w��}�&����U��tO�~��F�\� �r
oY@3���Ϙ/g\���3�>�9Ǭ�΁�[�s��`꓿��ld*ŽrOӛ�#٤(;��|�r��L����~YN���Fi���<��7�V�'�J&������|����Cr#>�=���ug��������}/�J�����Q��r�
��5٨�����/���$���+NA�k�c�)�w�Q�},YrWs��6�Aj���Y�ع��-�WP�{
�_��pO�J�4����O	:KO��ϟ�t���2�l5���hT���S_� � B���%ت](��$��R,oſ!��VfN�7�����F�m�F���.��g�T�)� pJ݃�	��{p)�ES�� ����k$sP��Uz}]it���ܔ�Z�2�h��Q����׺j��D�I �в���Y!>P�=Q7�]���8�?OZt2�)�JQ�+ӿ�D>�_���W4�L��G,VЫ��*e��㗶WF�s�P��4j?�����:Ζ�H,;=dЖb�tZ�����gʗ_֕��f@P�Z(S`D���	�1z���	�%����(/{RUr_�L������6UQ5�)�S� s�߈�ҏw9�P_����]:�O�����sO9̝�8�3ú
����eո��/W��Q��eKl�	�}�.���s�~l֫�}��#�we�.#�HNqԙ��l+���LA��Kn��Z��xM7rJ-:�p���0��͜;�m+I��,�5�@��^'#W��?H��0Pwٚ��keV7#�����:`?\!y4	�.�[|����B+H�^b\ 羬�3ͣ���1�P�e�aŏrp�vXW����mL�[�Tܲ�~T�KB@��o��@���$}�# ?��A���G(Q^nG�
Vib\S؃!V����pv�ϓ��F�(Gę��y������Fp��C%�a�QD�[L|k�Ƒ܋�+�Z����[Y���I>��ڰ�!a�������$HgѬCf7ڈ!ytyo)�>��SA�F�'6�5Q�"�3&��hx�����ۺdQOhN$�t	�|���]%