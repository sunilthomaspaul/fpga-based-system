XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd������S_%�ì�6�kK�{���~[�u��Ds6��j5��! $�tO4�|�x��_Ih�����u���Y��Z��ܿz�s55��&N�sZ� �E��f�;!���S���B}v���5߄X��"5-���V &����=�S�7�T���!l6%�P�OƄ!��6e�V������UZa@;V��o*�eAs#f �J�~���<��#Ңj/���M�rh�`>�x=7>������PI�/��|���yn,����!��'���bT ��`���hK���1R��d��PdJ��`�԰�+��Q���g�hU��? �沌Q�uL�>��U*z���%��GsS�Tv�m��-�ިV7���ޑ�Ш6���"��j�*J���P�c)���=�H��X�%'�'@ުJ�|��X62�L�I](e��e�z������E�I �T
���6��3��/��,�JY�'�!�C���?mU;gD�1�M,fT��PkA$,�ކk�A^�BCY
���ˡ��-c��B��dFD蟺P`up>Y6T4��L���e����6��l!�TcQ��0��8��4:�2-��4��_��eoc����+��ʜ��X��5��C�l��%BRI��w����+��z6�B��	�څ/K��C���gm��Jʝ������^�ʋ��2�ï"���½T���NPO���^6/"S&�@MאNs�)�W�fz���f߾Yߠy�= "�e����F�g)��Y �Z��� }֩�XlxVHYEB    5571    1410���-�*i�Q�Š+����#���N�u	�����ڃ�ͺ�U�Uj�&���Y�(	gޘ*��{�5\����N2x�MN��?�_=]�q�r�A��
j����Iu���S\#]аWT�����U���Ι/�_��B�R���+3	ϖs�u��c�"R�[�	�%e��P(��"�D�D���Q~��?��f��m�6ݐ ���GC��@��
��-8�^~����5\��$��M�T����t���B�L���Z�4.�v�Se
إ.��6��y$hV%�[�d�i���9�� ��6S��K�\��lՕa�֧u�u�N�o��}������
6)�oOI�K�M�~=�y����(��K���As�(�Q���]Ů1�^��`���A�(p�]]hl����Z��833� �!�'X en�N�,���W3��b4-T?ަc��P�V�~rk^W���[t.Z�{�V,��4y
���[$� ���H:ɴ�Y��r\E�Z�A9�����~���T'��`Z�H���@�)2�S��o`��KBҗM[Z4x��Y�ޭ祻<8W����B�`�_�_hEK+UG܍��z��ooz�]q["����f��R6Y�p9�p���5Lv�	�D����bA'FZ��%91� ��m�g
3M�8��Ia韁��
tE�^���x@N�S�W �\M|�
����阇��	!ϱ��'��7�.@���"L[x��NJ&fz1��8GH�8����C�i� ?���K˅�-a9��n�?�3)�t���(�k7Ux��i8���Uyk�K�����ie�	��q��l}�f��s�����ЈJ���������)���ࢸ�N�@�i�>4�G`�J�d���H���g#ڮHwam���~|攡7��߆����U��.����p����`�Y�C���'� ڥD\�~1�H>=4��;���d._?�t��m�h"�	�υ�Kge�j�y���~�P�-z����v����$�d�#��j�l�m��J��c��5�H��)C�sP���g�н��6����=����S�״n�О:�6Mj>u�W�9y���w�d������潫�ж<���-͏��ř��yգ��`9���rWs�NՐ� �"����P���n3�=N4A��iO�)��t�|F����w�]����3��s��X6쟉��V���x�;��R�>b�O[nI��)���
���zwhL�a�#�gZ�([�h1Z��'[M,��oqÞzP B�e���ȼ�/�{$�g&������^10D����۠�B"8�+��|d:q���:������47*FV@3j2���d�w,
�p�����}���8�$ B��X]E,m��*�.>��R���=1e?[+I|��g�s.ش��}߸�{�`���Z궮�$,��i� ��^��q�%�6M�F;��H��M*-]q������fC�V�?�������J�U>l[�Ϧˬ;X8i��������"��\�n� O)�:|kU{�_�Sȳ�I���\�ve�ԫ9��&�x	mf��>ok~�������6s��h��(U|ŷ��,�H���;��h^C�є�A��!!�:A��f<P�G�츲Vd.4?b��X�n��b�Nݹ����M��w%Yg7jJ�ʦ�{� j?*Ut�ᕣ��?N�lX��)�}-��3v�i%���׎2D�AM�Q$Z�2�}ʡ�d�@��uet$���ҥO�5��Q�5�0�?��R�^0��a���Ba6|�R����n��'����`1�@� @V /5�⺔�Y�o�08�~M���W8^�d��U�	��ň^���)O;�Ԓ�E���b�D/a�~؃>'ڈ��@7,�R���@�-�;��;qs*&Eɯl�"�N�A$�ô-�]��2,��)<"Im�}�[��4�	r��������G�Y��5���5:���c-��W<�7���T��a!�#�&�~��ip*M��
�BE�M>�ٻ��!�T02�W�@8J;GO ���}����y�Y7��k�y�_mY$�
����ulO�_����?��~�s�o���׫2ؼ�䰞.�	�w��r=��47	�;̽c��#�4I�߃^Wt��)�;��չ�ðO�c�u��L�5�$��d�ͬ"���?��?�p~�P�MĜ;�\U�֝A�-H��a�8=5Ʀ��Ei��d�����I�����U�w���^�i��Ӂ��٥�o��b��.�H��������W��EM+y%3���G\�`��B�h���V�Z
y�6o1���Q-�W��Y��.H�xw ^� ��m1���7ӕ#M�ZK]�$1,NpF�����Xϯl��?Gv�" ��s.�s���*=��w�R��!�"��5�Ֆ�*���ޯ�F6�: ��蒎wG�p����T��� &����ix��(�d�GOrN�+���\LW5��J���J��=��j�4�b��^�i&(x�l��4D�����rg:�}Mb��|@�����ڿ�9���3"��|E���2-S�Nޗ؄�6�ׇ���5�9��S��r�A��$_3<W�0����]����K� �sn���7ER���)��� �[3�  F����σم�c(*Jg1p�
�����a�Ѡ�7T	:}.���	�b?X�|!���#5L�(��ҥqϑ��Fc��)���uT�1;��������%2����1N{3����YĆ��)%K(�sE�h""�n�F^6�B�x�� �m��P�-���<,F�O�gpت&nv>�������:���!���mG�k�-��Suߧ7�v�"���O���a!͕�b:z�'A�<P��b��3A�=���7�#�7�@�g5���Hh���͛Ժ�j��R�����KOb���P�g��9���Uɐ3�@�,p�Q���.^|�;�s�<l����E�u�؇�6Zz�����
7E��lvo���k��of����((������v�-�"��b�Kjg�#���Ù.�O1���@�d������G�XB���Ǜ<�����X?�<��je��1I�L_ؑ�p�;|�;�8n�D��-.�M��	�`$�G+��\���.�ș����N�(c<O���c���?�ۯ;O=���Լ�e/���(,�)&>T�`�!���z�g��*o%�2�!ꩄY��a�p�i����ɌbJ�ܿ=����Mr�=%Zd��I{�"Α�x��z�]wÁ3+��6�W�	$+E�X�[�Â,J��&��q��&_��D�uK�ڮ�:�߶Q���YPR��K��
�]Ɵ���:�)ވ�72���A��\�;�>zN7\�Xr�t��N��m��ϗ�B>Te�������~���NPc.�e�Fvq�����o�;���KZ8Ό�j@i+����T�:�)�ѸC�]����G`�.������^�<� ]�@t�}��V���H���hj��n� �&��C�&S�,�R\z�*�sjN[�1��ݡ��%6-��|��hC����.�ظ�+�~�����Y�xF2�M;H(��$v9���� dRr��2�>�W��{���n���eĬ:�ph��eR;TyT���2u�{Q6�GK�^�9J�C~LT�aF�`pw���^ʥ��ʦ��%���.//f7�'W<��6�}�;L{v��N|��`�u�Ȼ�8Ԇ��`ׂ��p"񤶐Bv@�Ad#?">�̅IbE@�*�D��lKoM�Y~ܱ>��~���\+�� @�E��U퓫�M+�Sl�9����N�(��YX��(�WeIbg<96�*xK�Sڗ_�.8��t��NU�UFV�D�lާ��}7*�R�1ɠ:I�_�2����98 �>���� 0M����|�S��������VPw�N�#߀_� ���A�{;��~am�/ڿ��E�*�ȭ�smt�BE������~�J<��_ϵ(HfN C߲4^�F���M����Dxև��(�Ec�{��i֞l��aX$qX �W�œ�N�i񉉋���^��V��ieT����� -Qu�F�C�H���o
[)t ��xp��f��i$�uw����r���P�U]
���?�KY7�c�/K�]�fX��.�`�-��_��ͤ��mtm��2�B� �� 9�,T`5���h�Dn�kE�~3����SGG�V�<$3�b��WX,%@�N�{N��e�s�;Fv	��pȽ�lg8<&�.�9���Aض.I^�ϻ��CZz���WV�IC�x{6?N-M��.٤U�Ɗ�{��8¿19]Lz�P�E5�>�Z�2nFJh4�Sԭ� �a���7��>�㠲l|����mί�Ѹ��D�nM'���/�H���z��/��f��=Y�֮�;����k>H�ІJWb-��]w�a��P� F��(ٖlqR��
�P�%����w�Tq���Hoy�w�w�vm,���PD��؃�iY�:�M�,�It�u��+ֺ��r6��3�j�#(��9n|�9�V�Ӗ"=���������N�	���	�X>�WS��Q:��o  �5���T�s���4�++�}���̾ڙ*e����/�q���ի��%7� F���B2�$��}*���-�VǼқ�6㩒���Bo6+*~u�|d'Ktkr菲we��JA�	5�s�;oK�k��� �1�.�
_נ����q0w'��iߥ���6��㮽�S�
Y;�X�?k�o�o�W�*�J�j~�\��xO����ݱ��7�%�q�_��S�Ļ�T`>>B�R��W�h]��lT��d;{�1�~������5%Ru XC7�q����ymL	�<����y&+�����z-�c��v���CM�ty�3��:+���/��рW�!	�œcx��_A���y����|F���G=a$x��=WUê7�.e^�a‭�lx�z� ��1�;��3��\�w{�;�x����;�4�<D��U�AO�C���6��x