XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���=��Р�מF�<�tz�I�����[��J�S�0�h�$H�B�u�j���S�� X�O�l�s��G�N����4ɒ��5��Y�]\36����
��D�^i芦���m���[�ǌm�z�C"B��`B��a�8m�z�œD�����B>�#,�b�S
;Z3��q%�¶O�"��T	R��@�^�|@��V=���2�њh'������/�,:sė�aunwz3��5���oi�_�����6�$�������MGu�ϻp�Xm��q�IKt�P�D絝��U���Om�qؽ��ƢB��]Y_�!��>ϞC5�0�@9�B�9R,��c+t���o��g�,���MҀkhmX�+g����S�'�k���J�K`�gN��q���x�1Fo� o�%`!۪�e]��;�l�_�h�=��̱�$�UgÜQNY��W܎|R�?\Q�M�9�G�p�;]�Rȡǽ>4{JHN_��������zt������,���縮�I�n�"~�Հ!�4{@��V���ҎLV�HFFW�+��ۍ���2_�����P��)�0��S�V�z%��x�4 u�V�B{����;��!�c��c��\�r@��Yo�q!��!ޝ�;���զ�Ե�/�q�c*;�e�u{G'`�^����������J�}� $A�QNȥ�t�qX��Cѿ�����kר��6DK�h�CYck�=OKF���O�G^�@�z�}�2.QВ%�'�q��P���.�H'�!ll7�XlxVHYEB    bc57    27e0π /坵]����9���Ì�y⏕ay�1΀���p��?�_J��^e�`��{�{��۞kӣ2�b1��T����� �'	7ΩV\�v�_���ߘ�G�%�x{���fg� �C���3��Ŏ�W6�,3�鹃�/���
<�aԊ1e'{L���d�)�֟[�</�ĲK:��HҜ^!"�8�򜳵o�mMI�%8��I��g��t.�)I=p�N� � /yg���`��9�r�m���RE���T�	��Ob�Zf�VTμY�����,t2G�+�ЦU��|���!+α��:l����u��C&G�,H�pٳ�
F.�HvX'�s[�)mԻ�!H�� �l�w������P"־�t���Z��de�>���E���hz�ܢ�r�#!����5.H���B���	�����UyX=P�����߃�{ ܔ���s������U��GS���G"g���}o$}������������ÿ�u1�
}0�͊%�?l*�9�Y��~�/։�c����մ��R�s�1ǅ��/��(
4H5��dN4˗��u.R:R���0�D2���j��`bkv�aNAY
x����r�<�hGV�a<1y���u�J�X<K263��N׋�W�a����9W�X|"]��_`|�N��?	���b����|��p�J��%�+1��z���u������1烎cPiw3�tmk�8j�n�v�D�YX��d���s(�;�^T�?��-�%\Q�s��CE;dN&ש��z7��@�H�v�ͩ�:Bw�����f��l� C�N=]��{=��F�#����o�`Ͷ������6�Oy����ӫ��|R�F�uS^�ӹW�Vo�	z;K���tJ��v]�>�9>X�]l"�bUչ�^���T�>��z=H�5ǇsΉ�J�Eъ��bX�-9)30����a	ʏm�U'<I�(�当{�G�u�C,]o8�4Vo��X7�#�����m7�~іPެ��Ǆ.ci�tX3�-���#�~�Q��Ѧj�: A��Gd<i�b�g���r�g���������]Yb��m����,��FN7-O*�N�����ZC6&�Ԍ�Y�N�:���I�æ�<!�Ñ���0���N�x��U�X�����Wi%���yr�2c�[�_5��Gv7?���3�Y��k'��y���s~"��S������qp�%~�6�����V�����2ˮ��H���1m�*c�K:^�bv�e>��@�Wuu����Ӥ�5�.)��TL���QD���6�9Ș��͍ �-Z���=#o��ܾ2���f���i����rj��d�U_.�gi1E�2��c`䟟D,�l���	�M��vC~,L�	�,y�b�]��_�7Xny��1�}P�ϟ�]A��5��E�,���Qs�G|�kz�!�2U��+/�i���}�b�p5�r������Ȅ �^�ac2�g�:� p#�����A�t�	�rB������r]�n�%I��f$#2��������Kg1��X��_Zq�J=�
A
�XEGw�\(^����CC�m�^�^W!:^��1���	�{���3�Ǿ_���m!a=���� UQBq��T�l��h������ij=?���7T�$��5E��t]�D���#�8�Z��67G�rX�m� {�:�f��hL�۠�Ѐc����_o'��A�.ʼ��)c1��^���to���]�zF��[g8�vg�<䵕w�AGGWv-}�ݮ�'�x��nV<L5ڍ97U����x�J1K[��d��l���BN��iGB�Q� NMz�4Q5յ��/���y{´��3�AѾ�����E�g����}<��Mt��*Z��r�;�l�������u� �����O�h[H���-�,t�;˘�[pOT�����	�TQ��ʯX%Y�%�>1����)&�����.ĝ��[����:Ǿ��
���F�ఫ"�	(�d�]im�q&� =��y����`��D0��S/�
5���2ݾX'��3��Ʋ���;&ϙ�������H����f��j�x�
'^ʧ���A�5}D��*�x�a:����x��8E�)�J�@���c�����b��x:��MP�=d�t��1iһ{�b�R.$��/\�[��Ԥr����%h҆� �4d��L��.Rb$߽%!Q>�A���?H0@�K&��V�c�"dv8�����le'�I5��׵F�H�VH��Y�Èe;j*��P��}O�Oh�7�`�h5F��eF������g�D�l�%Q⊟?���O�㟩y���tjF�����2	ͺ��C��l�J��1N��Q�pa��G��K5�ِ<�����&���ڲ���y6i-)v�G8�Nܢ�:\tP���kw��0ټ����˲	bwٗ��0&L/j����|$/K夓�����JTزZ	r�VaPP����E�$�F30]y}��Ⱝ_���H��ʿ�$�m�O�?��k��8_ۦ+[E�j����J�i�(��)_��'HL��qO/)	\~(���p�fL	x�)h�'�;��*ݿ%h���
qSB�`����4�v�%��R�^7�H0q=�P�£�
>P�IK6�jٮ8"<�U�� �ogx�}g��]�JK$��F/����_�� ��>���!,�%�R7Q�y�p%�H�u�à
:�5���#�^���2>���}Phsw�8��ŶH���mi��G��hj�H(	��C7)��`2��?��[ߖ����Ro=^� �d�㷁�ã�o�^��m��Σ��v���ܽ�[���,"�ҹl9��]{�}(k��b���a����tCzx@DZ�91G�<�?j���@��Xoeޕ�g��o�e�$&Ă�>�Yq��K��!���qW�`\u^��������wMj40�M5��{R�:<������C��2�_�u�޽`���)9�?m?�9�<��/PN��Y�AO���r�{�0�A�+F������L�EXW�
� 1��_C�V�#	C!��\�m�<|ql���ܮ�����G�2�����c|���`��-��q��y���/�1���%͵v�$��k��>���b��q+6��lA�U������]+d�{x�i���V[�:��c_>�d����/�
2RᅉL�����);ġ�3��/�5�ccf�	��49�4:Ʀ=ݤ�&��e�8a�UU���p��[�E��1%!�n����Jp������SMz�I���;{p�9�rҕ*�j�5�\#���D���ݪ\u��@��c�S���E�w��߁r`:�\@��N}�hBf�a�q�!Gf�{�r8��y~�+�῕�}X憩��<rt�<�v=�K �<�AYfh��F��ʠkYbMµ$��f��{�r�o��}�Ic�ȇv��Gw����G�����^>8v,��	��\�׆���@�z��z/�{�a��h^L#�t��	<+/�h��L`�\)0��������u$@��ة��&��\�}��\<����N�Ih{q�;r��~���F^�-K���dV�_=�Lsg��G�%{(�xô7G�|���R�8���]ǄdI5YK�A�A�;oy6��iqe�itK���W�Y����6�¥;�͙�*��l��k��ךV	� �c��*)�No�����0�����36��2#U9�}];H��I����ܡ9�)i}�m� ,'Rr��������Qtռ�+J|���fyYg�Y6s$D��u�-��ACؑ�Ϗγ�8�	������O��İ���"nHZJ� ���k��!����	U� O�����g�K-�>�a�����	��y,\7ʹ�<�G�zme�p���#GS�i�;��g���u�? d��qd����Pؐs�Kn�E
����d�4�u�z)��Oaq��yӾ�����_b�K���d�2n���8�r���|�&�a�Sa1+�GT�PM��e���QN�x �X�蒺t�b9���|�9c���A`����s@y�t�l�J�渿��������3����m��!�ARxI1�)#Rd�d�u;s��7:�����
�g�G�Տ���'�H�{J��1y��x-YҊ�SiQ�o�-�_p��F���:�&h�-���|z9���C�$5]Dc����Oa"ܡ �9�0�{~3>���:$l�#;�,-�<J$�,�tq$���wa�6��k�b��T��a1Q=��Po�M%+$�I�� I� ��$rb�??w�%iߥQ�q_�ס�m�`����ç5d	.\t��Z�@8���ю��NBQjeP�eҨ��w{�=pM�E��vҭPu�0�{�OdC�E�<VN��$� #x�+
��pZ�c��#7⢙����7x�^�͞Ì��j{ysc��8&X�[<{JSPP���`S`��#K�� ��M�̐u_k璉���&������'��LM�����v����qt;\��ǥ@�P��i�E��?5�v����ǹ��� �m�;��9�=���H+�ߕ��߭��1�m���2�HM��sᕢ��A-�-���`w��j�*�<^�������WE�����/!_�rr��EeC�8}oh�ÃUI?�v�����HpP�7!���PnN�|�.���$���H������_l�r�D���6 �](E�Y����
u��gY��{P+��e�>G��+�15�-/SS�/�k>���i�8��E[�B�������e��@�M<a)�&^	!e���<	ysP�3 ��C{f�sg�������1KS�O�F�U+��&�[��	P}As����\-�C{<��� �׮e�e ~����6��ϒO#�XD�c�׾�a�5W�$u��R�~�߭ ���\^r�h��͐W�/X�� v8�7�n�Փ���L8�Y�[V�$��		�B�����5\W`]��*�ٲK�q���^�J�w��C�oH������AC~yw)wq�1"�ϩ��q�m]B�	�h�-]TV5ȓ���+(od{��C0$�%# 	xN�Q�fCXz8�0��#�{4�ɚ���J>���;����H���QBl�_<������x`h��<�`�<y�u�������C�u�@�_��eѤ ��.)ɲ0���l�S��	¶�#�gy���~f���������P]���2exi��T�4�}��Y=�hi*�x}��F�. z�������!�RPX�����]��v�/z2"�	�H��뾰��2F�~�i_=���B�E��e?�%��e�$��/E��@͝$�:��0�d˲�o�ZuM���x(�d����Pǳ T�1�9��R�}��^Q �//i�*������%E��of2��OS	4��ڍ��%o��n��'ͣj��M~/ �n�M��Y��:����� "�Y��l�-�E6��{�X9�[Iʎ�<tµ��Q�����y��7K�^b*�)�D�-��ઈ�݄�e��1��ijE���e��]J5���^r�{|�,��d�i��[z��f-��\cýޥÞ?��:'���t5W	����6��$J�XZ8X�L�D�xdO�fr�P���7��\>L����&1^��,� �����0\��1���	�O[��g�H� Nc/�����4����Fy�ט�����W��4C���\�]N�A���!.����DR��5�:,0C��x�&�I[���H�N.B���u��a=r�A�K/�h��)
#i8������l��jA�ƕ��N��8���"��^��^hK����%��,��	�c/<�(kL��t�9Mz�����]RM�ɚ
���j2�w����ώSɼ�l@Y�g�3�gZh]�O���f?��DEB��q�yv�\b��*%J��I�P���?b�".�����F��ŧ���hʥfl^�$���R���=ӿS�Te@��Q�y$��u���(hU݊�9q�Ӎ�@�ٗ��.��h�Ől�3Rbr����y��4]�ԙ�;{_̫R:�3&���ֺ�ΓN?җ뒶m��5�N�̠�6�2�4�/45T�-R���:���";4:	�v�7��:^��mv����w>�D�O0�$�G�� 6��e���h�ye�R�,GX��')�������.DZ�����1+��oM9(�IxB�ۯ�҂�k e�,��Y�/z��,9T��Q��j&o��/�޴��	���TE6�8BD��%������Bt.�1�8���ع�G�o1��@���m�$��C@�]� q/��ͼ�������f���mq9D$-�}����>��,����c�.�(��"�趉��MoVµ0����r4��u!D�\2Ok��x7�@�ncOY�'<м�"��~+)�4��ӯ�OB&�kf\���|~T:52^�}��ˑ�{�߾(�G`��F�E��/�Ģ���v�w4�g�$�k�=X���)[���S��������ф���/PC���p��_#J��8?O�8U$�W_�ϱ�>���t�Tb�N�z��f�n3ؠÈ�l$��L<p1$�]P?�hI^VR����H���g;�A+(���ճ����`6�>:kL��"�$ĺG2J�D���11w�u/Ì���R�8�䱊���vsy}D�i��f��nBe���Pz�i��| {N��x���Z���f��]Q��0βW�����7��$�!7�syM	Sv��(�C���F�
�b
$�!��7�m�ZY��;�m��PAl2Zٱdi��"[i�>�i���_��+�:,`�W[�[%b�_оfo,m�u�(���z�Sٔϭ��9x6�)����U�Ϋ�9��{��}�z�:}��v�[W-�Zj-1g�����h-��wa�g,[�1�:EV� �k�.o���N}��I�&u��Ϫ]��8�_0����K= m�?#��6�*'��a]��)\�ce�Qw�4�6����-��46������3�Q�?n�g`��}$�5�c�r㔍��L~�������n�s;S�e���B�k&�^r��I��t�D��/��E��-���aPr�D�����n�Q���9xg'�,`���h־���:>��X�
9�߱֝�21�0~t�����f�Q�I�Z�M��[�W�y[�j�G�=��&x\zG;�h%Hl�0�T�F�g>m��X�/Υ�,�V\zn���ȡ�׭�w����]�S�Ez}��K����m}��dǄ���{��J�إr�܎���=ˬ'�`0V}@f����js�Ɇ�蠹 ��{%�B'A�]T�+,�f�@d�<�QT��D>[�?ܜބ��;0��F���ct}c���3R���Q;W/��6/�r7�b��t�jN������94�)}J�o�K��T���r�z	���xa��7:'��j��3F�J��&uC�v�fєA����[G ���jk��ޮU����t��������T��l8�������/
G[8퍳JÍ�5,�eV�"��+����7����>�u���v�,j�� l	$I���)��0lҲо���B���5"�B�j�}��+������;
�/(���|�_�������� '�meq?��>�n���FVi<�����_-Q.�T!�7�z4F3MD�W�'��1$�I:0H�����J-cTM9�Bdz</�f�QM�ⵗM���&ܯ���vb��꿾2�`�����)�yӓ��j������L�6�����L��Bbh�c���G��#��
�ɪ���� E�$|ѥ��yB�h�10�=��[L�Y�ꓰ}�)���fƍ��"L�%��'ڎ�څ�$Aˆ1 ������15���{��%��^��A��L�[����QTs����yܐ�,��/#< 7C�14�P5D�7��ƽ���^.�	�Z.�*v���ke��J����>�M�L��Oc�Jx ��,�H��#�`�_���xP0��*\:��o��aC������r}o`�7mFy�L��cN`x&�=<�db�6��ɮ�_>u_�۹�;�Z4D�Kj��{ǆ���B*��+����hф$[?8[vN-�+k���k�O�^����Cr�h���Ã�s48��ͧzǚ�!
ǻ(�Ԃ��o6Z�	��~2��o��ʤ��5 �,��'�'�f�(��-���"HUU���rN�6*SV�b��6ɠ	�� H̢^�qb]$1.�(���� �|�q/_%.��	d}
�޻P�Sր��۹^a��;�D�� ���;�aXd�$\����3��(��1�F9�"y+�Vz�am��c�Z*7ϗ��_�ϊ��Њ�I�G���<�0�;�\w:����]	f=AO{X���B��5��o��~m�eq�{/�5D�`&E�����i��?PY�����2f�	_�ڪ�Ğ�?�g����)`k�!��!���*RC�Ὄ�a���[�Ep��d���Y����8���p�eeѡւ��uf>;�K��wv���s��eH��燅�Єǵ:��Sނ�����ә�S�M�]�K�!E�~���AU��?�<��d��
�/�*��W�r�tt�t-͒�A�9iCN�'�	0}�@Qfz�F8�ez��2��l��݄�}�̝�!DT�*[�b݁�F��٭�!?�hѾR1Z�$��\ D��T���q	�
ʓIM���q�Ek����ʋ�Q��c�Ể�z��D�r�R�¢�Ȣ;n�EmU�aC����gR��5iܢ���$�/\~��\n�aʞ\a�����R���#��75�JK�A�;}Y����-��7ē��W��'��>��;�ͼ��K�_��=��TD;��:h�#�&�j��|�L�|U�&[�Y�:���߂��k�,5�Rk�G�#��͛S�T�h�O�ɦ�
�̙��6����m\��_������wW��W��[�����@PG��#�;��A�� {V���a�4�r��' �����'z��,U].%T��]u�M5���ezӇ�*C��1{Ӛ�NJ���I�B��Wa�������j�~��آ7 Wۿ.k������
�&K��~x-3��7�|a�`���*b���Z5���ke�M{���b�AN�:*�=t�
����F,]|A&ԇɤb3Ep�o�����"�T�ʂ�Hܩd�����@�7��IZ+1Z��уՖ��-�%�Q�X��y�Y�Ý�*r!n���������I����=�K���q���E��x�*A�,�6�kߵmwX�4������K�u�?�,&qH��p��˴���-�-F\fYgQ{I�� >��n��YC��U$Γە����WA���,^2�³W�*&G&I'_��WL�U�ٮ�,�r���}���n��<��p��6b�ňB/)�a�M�Q�o���nj�p+�b�B�qX�?��D�k�đ�6ک@^_@c�2,� ]���8M��k����`T����U>��YV���@����;�tj�6l ���Е�Xk'�pP �[�*��i<�\~>�mC�߿�/o�g�����5�n�UG����C��W*�B��k�}�~͞�hI~����fj�T����4dQ�����+i)w9@��{�k�6c��-�'d��>e�qtFǙS���(M���׻%�	�Tɛ{�[Ѫ�J-�}Is��׭)�T����=��1��s��Q?Ml?]f[��p�3�b��iP��t�6k�,�@��c6�푥"�#�V����K���d�C>Lߎ�����������5���OJ��t����`�DV�[]�7�V]��N�\���'�Tb��	u�kR�����
%�;���'�s�B]k�%[��"���S+���0�N"�+�2TS�������uK�P���~jZ�T4�̿��6.T�r��2�Q�h�`�q?@%��7�S�v���mF�������1�0��~6
��=�^ã��"FQP�
�:����Ý�'�N�G�#��e�