XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����H�inRU��?�(⵲�7W�NvSI�x��\(C���(�u/�P��.� NѪ�7���?�����Riζ����x"�<){�^�����Eje1�=�� �yAu��&yiA)}'Y��L��n^���)�$�
����=�E�<M����u��&������C�1&��i�����!ҚBO���vޭoo�]�d�Č[8����?���s���hF^�]�Ʃ���C1�<�9}G;�픨[1c��"��z>��9Yc+�^WV5?5�baFĭl�hY���A����3�b�χۃ�}5�S{J�D��x�naU���4�s�SF"i��!�
9\�M�uL�k)�*��qe�"(x ��R�41C�7�/��ƖܽS���Jcb���S���X�{6��=��6hn��P8������ݦ��}Yϧm�e�&������zJw?��X0��x�X0��{.��=��$��Z;�%�PCO�vk��4�v�S=�.�Z-js�q�Qv��@�8�KL�^�����$B~`�)�3T�N��K$���.��q���#��~��w[�������dx���7�M�� �c�U����I����B׎{�J�GGqŀ#U�Ӽ�Tѫ��Z�J[:�>"�B ہ>�C�N�\��~"�ӱ���.�o3NZ��g�qqQ��U'w	��6*]Ps��(���;N�������#���h�&Х�UO;��[�3����
d��g]	5��&;�#��"{p\n�[��Q}9�_�[���XlxVHYEB    203f     a60]��� 8W�Pݦ��S��FV����������"��-8�
fk%Pŷ����A;�`�ȘC�{�ݜ�z�����*P� �0{#����,lgn�@���F���)G�Y���z�)�_��s XP�Y�*���^'�St'r�+������Ș3��_�����{C��D�Lk��%>�\��A���h���/ ��s��D�,��Xwx͓�}(�D��>�{TZ�d��M�C� �E�8��0� ��t���|#~��[� ���ݼ�-*���:���⦴�QE�V�1A���Vs:��I��J�v�������'Z��C�J ^L[ꔇ�K2���� �b������ڟK���/�1Q!�
p9�YI�2/���3Ns�C�Qx��D��L��6�ᆸ�dv)��	g���7�~�O'�7�N�:�<4'��FZ�I��j?.��� �K��L���Q��G8~GB���sY�r�1�I���C�fն�rU����;���h�*��/���,UG�BzM�O<�f�n�9'�w�qL����B�m(q=)��}pϐ��Q�w4��-��<O�&	#�无&�	zfj����iL�d�
&�����-Q� �����F����RbH:�0q�Q�'��1ܹ@��iE�`��;M�wb���%�[ �x���gg��=j?�ƛئ-kBŨXt�.��ZƗ���0u��9ߛveP3�R�op��pC$�Q�&�<��j����̼��v?.�w\���^�8E�-̕fT��|�Z{�V������0-�I�f�ց�Ed�eO2&+N-պ&�0mJRnJī�R���e�q�$i�'#�6.�Şn��g w(���@�*W�~���$}�+kw�S!J1Q�����]�����Py�9�؞��s�JñDiOJ}���3�x�r���R+鴶��&.������h�8E�_�H;~4_Z\��1Zk���8��C�(���#��:�PrD�gb�$�j��Z�-�Ȇ�>N�-��k�p��/�XR� �����L';�熑e˕M�9�� `�����R�d��)
9�}��Jz��޷��X!$����� �s�X;�-�����EC� jm����)�bf�(\��qFT�h��J�J�Ĺ4�i^	���F�Z8����R"Y��(��K�Ɇ����e��$�#塙̯�F���/]_&p3�uo�]m��;<`g���r�>�Eq0��&p�I�-�"��"����rk�8^�@��"���:M��O��α�'�RUɧ�)��zd�t��ڸ���ū��Έ�$�Hݲ�`(#�2BWV��ϲ*�~�"'�l�q���x�1~�۹�on=ߞ��c�ϳ�1X��h"&��*ZZB��<��I��5Dy_�˩W��L�w����|��o�S�vϹ�^��j�D�~�@�"��d�@��:��a�pM�۳$��<J
�s�[����}���F$�m�HHI�' �D�9D��zӸHq��Md���vI)r��mI��~0�!�����m�~-����S�5Φ�Ƽ��r�a�R���Bp�[iĆN�uCf��I���;)b�3�I-׵G+�ʭ�&�S��</?�k�̅��^���cW!�'7|���K	X�������[���b��H��,pdR�y�LNG�
�uԳ��	���=����.W����*VE�:�ܘ/>�Ʌ�jt�<X$�����P�J��W�Q�vx �q��4��v���D%�:��LΞ�<`$�]N��hY%�������ˑo�3����xA���R-߭�e�b�H|N��g-����bg�ܜ���,�_���DS���Ze�}т��z�x�"7�bә��K>��!ێ�~^C<�l�K_��0���(��t���@=S���mv�B^��pdCSj����B��Y�6A�b+������i�C���]�|i���o�,���u�{�ԔO�*�')�	jt�W@O��{�T�1�U�
{�t[��f�r�����To�Q�Z�+wε�SR�1'���~��6�Ya�@8�^r�*B� ;W��Ir������i"	-��56��Ҩ%w�������50u��VE�"1�W2�Y�m-�ˬ��C�k��a��^;�\{�CG f�23�l��[żTO���|����c�_Rl�lV��'n	:M-��N3,L+�5@�s��ܤt`�����/�3�3���VNM��s"L"A�F��v��^?'���o�[I��Z�.��)�8��H���H�Z����U%���1v�믺�Σ%� Rny%��y�_��5x1��B��$0�떘��W�)�����x�g�f7`�m1�5Wܣ���FHn���G6�m#6��
<�9�EGfְ6Eo�EZ�x�o$��G:S�zɷG>oaѴ�Ĉ!��Wm�Jxd���Gg�/�>H�N�noѲZ�G�np�Je���ز�\*D�b����f��tDQx�A7����9J.L|�+zU�|PEx���ªY|��nܷ$�=�B���)KQq�R2�������-n�
ٶ�,�������2#U9ʯ2���G1���a�����.�x���w���DU��'��x���Oj/�˟r��&�O���