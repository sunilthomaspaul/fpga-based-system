XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��(z��Pbw�D:��*�o��5}ϴ���d�k�l��h�쟋�5j�ob�>}��%lB��C����n�Ǝ�U�o�����X��-��ԓ�������.�#VyM:�
�k�D+�M룓���ݧ�;L5���������ԃ~�h <�݂x�pҧ$b��j���)L;�Ҷ��p{�61��)�t�B�Q?9�ԹD�P�pht�Q2�*E����t����'+2Bs8G�F9���P�3�_`m�v������n���U�ٿ�0�-r��as]P�Q=-`�?|.�R}�9Z}�p�wqkL�u.р���v�ɖ���E|)P}�h?I|VI�5����H}̘�21��_9�K�J�t���h5:�^b�{]���7�v
�������Q��}Z5������!~�~ ��t�i���M_� R|�P�S�`Q+�����V2��ߩ$?���8�5CXP\���F|4�3��W]�1�7�. Q��wZ���>CP�Q��,D�Kr*��qb�=��+?�����z���F<�?��'T�{��kI�0i��-�i�����\�������x�F�l�!:�)��4D��
 f���D�e������đl�:BQ�M�D7�#^����x��F��-��\��#�2B>�}v��-�g)ڼu'U�Vl�E-jґAr$5��wT��E���Pߏzm�" -��� X���:��HVr(�zs����l�f�l���A'�fw��h�Eu�do�ܣ@Se���Т8'��:0XlxVHYEB    19c6     900�{u��ﮫOgK�f:�Ue�0��zH�9U�8ǻ�G�MLux����):-q�����ӭ�g��s� ߏ�[��{���ps�*���A�zuP�A��VRc��������=ƾ�ˆ���~%C�vv��&�V�wk�,M��7�P�Q%�~ݽ�9���|�J�1���Ѥ�D���������=��s}�y [�sV?�ݲ4�h����(FI-��p��}�ON�4��Ӥ��)1A���Т��U�3ۄ�/��;w"#�R�����p��oz6N.2l�2�ʿ>��$?�E~(�CA�fP�ʆ.�k��̩��eKI^�p��O��d�pc�:C	2�'"��Z��w�4�9��n�p6e6��Ce��0��]K����J��=B:��>�W�˩B �4b�p�i�ܘ�Ȳ����ca�&n-���� �t��\���Ds���΁��l�B�O���cC�{���u���ʅA�����ۘ�Q
f�G,��5+��^�5 q,bu�`�I|�)���=_�A�������� 0w~ j̔d�����e�]���_.���Y�O��ړ�S��~}�?�q��[��̵VX�k�h񄽶�VOg�s8TMS�=��
c_�M�%n�`W�l�ԙ�qT�[����Y ��M{z��zO$� ����}�)�K�����G�Gy�g�\�S�:�&PJ�MP����EN�>�ƀ\h�T����@frh�FņB����9JQ��V:��a��wO�W�6��'[�Z�����7>�f�A��E�Q��X�Z��Q�it����1���k���\"��s��z��q��j4�����҉���nd�	�1R�^8�x�?��SK���Qq;7�z{�<ru��Tu�A�R�x~I���'��w�Se�Zǰ�G�E��K[@��q�Y��'�nF�:�T�����׹2�c@�2��h	zʉBT�%�Y⇼�e�����rQI2���6�)�NyD��Y)�/�aȋf.�}��WFn��,��R<ժ4U?IQe�ҹ�)��V�K��`�I��vTuo�^ci��9M����Z	l%�.x�i�Q ��Uq������f/�CߝZT�݋؟�va��W����h7�?U���g��)ho�.랞y�v״IK�u�����pL�̠G����cu^�~����)Y�������!�h��(k�3ܥ�r9��)� ����y�}��@^Y�ϖ�F!�:�8Q�2P��4]~�լW���|ڳ������A�%�+�I���b�F��i��\4��ϊI-����M]�8�a���>|9�2����1dS����9ƴ��zCw�(�Z1UAvL�Wa�AIG2�Mh:�­��_�B֮��8-���x9O����2RZHv
i.j�b�%��{ׯJx�pb�^�
c�8���P�z�uP�RϜFa��~�	׭v|�2�]����ڙ��ZXV|{��um�!0e�����Au�
��)<᱔n��	{D�����t�����A�[Y���D v�x�[�_׺��M�^|x�a�W�����d�c��-/�R�Ѳ]Ώ-�������(�@���2�q�2d��W^QE~�����M�0a��5���ĴS�	F3qC猟��,��}�BAE_�o�|���d��g/J�nA�H����^�<8K�B�@R]�?�|I���Ќa�m۟G�PJ���s��H3-_���,E��c5
q�dn�� t/P� "��>)7W*̥A��Krݪ�w�ใ��8���Nθ��FJ`=��|��~��kcIB��m�|��d%5�K��V��_���ʰ���Rj���m+V��H'�({o�y�8�x�(|��u�uպ�Ck�K���!�wf�o
v�F��^�˷;�F�Gn��`V%	�����(Xp��b��6z��-��y/r1�"����ӳ6	��ުn�����i�0%��KZ������<���1�����J���Ta��N���~���pE*Z�0��E�L^��Я���2ͨ,��%O�B�ҕ�$I(=�<Qzm�w�l���ɝj�!�p4'	�O/^�u�{N%���4j��(�Z6�֛�[�Lf�;�`���Q�_����exd�C�1�(?� ���,����/�)����%[�Uw3�^���G����A� q��_��Y���\Hx˚��}��D�b�����r�̚��$z�M`gW�^�<_,���ϻO��3~e��L?�{� �ސѩS�C���	�F�s�U��"�R�л�F�sE�