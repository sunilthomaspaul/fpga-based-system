XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��y�(�n�c����ߪE��ζ^UM��x��@˿!em�6=�t��r܁��Y�ͻSL�q����6~ �;"�x�R��:�,���O>S�;��<y�Ew��o�����^!��\�a#�K���Hx��wh�o�鑸�(|{#-���[\7l��9Qu��j�ƺ�$	�f��ì��u%]7�J��1�`Y��o�,p��a�]'�1��,ґuM�<��J�*��͝`u���$=���@~����~���Ҕ)S �Ê=B��&|���4�yU�,?���{9��b���#:���g�d-�g�!�mx�: N=_�d0�cIJ{}Ֆ�'j(�靉�QDYFk�ܡW��F��ێ�'��T���i|6���ېY#�O�2������8��cR�*��ly5���j�)g��L���ۄ�_�wۢ�Iɴ$���1v�����YX�����l�Px߂�t��] 4[b�в�_tinU�*�_�N�_�zn(�#3M�v�ZǍ謺r���j7�y6�4H9S�"�/��~�d���-<�6����M�� ✜3���/Fc���g�ٹ��{�ɛKj��@�����*e���a ?/D�XS9#��>A��8�
���+�w�Xw*y����TP���R��)��B�zA�����6���2��Mؚ��M��S�݊چ�s J+�6��*��_����dZb��o5�����?�k+n���5�
��0B�w�p��pf��=�rb[.���Z�I�Hy�sa�R(��XlxVHYEB    118c     6d0;�A?����i�$Y�k��v�0��qg]���iŊ�;0�V#�:���C�M��N�+�Bz�9�ǒu�8�@��'XP��j�1���S���E�kƍ�.�����'�,Kݦͫ�\�{h�n��������	������x�R��.�6%��d^��ZTD w��Q�"��'v��%���zۈ�D$D�7�i*dD��9�ZY�9�D�f�E9��B�U���M���&�+4���
�z	��jŉ��K��0?��5N(\�V.����|ζ{P����N����^~����_<	��.��\���{��[�5�|�E]pkp�3s@�/�
fgܙ�z<P�� ��Il�l��㌺���i�9x��2
�G�R�i�$e� ��lL,��[u&�	<DQ�P�����m�d��1�=�4��l�X��� 4AJ�k�����Vmf8�g��ߨת�TNq3��Ŋ���g%�<�+���G�Q���1:�k![�.	�1��Q�%�?g�ƢoK7�� �*��q��c����(IǺ�'�mC	vΙd��(�s)Q�� 0l�5:z[�r ��?�L�^X��TŨ�	����ֆ� ��Y8z@���+@+~���O�hi��=KMŰ���~��b[�����e2 ZBl���z%��Ȕ���]����e���uԼ��M��m���wY"�S8��ɒ�� z�^˧P�)3�Ӓ05̿�s��CXd&���皴���y��ԬÆ. �2�N�"�2��� ��ez{�]iCш<BM�����νx,��2De�)(Ga(�$c�&�zeqK���v���?t޻�n�)#�����1�i�g�1��?�+B����:SdeggsUh:[����KlsJ����i���6� !���nL�:�����ny��ADyu�i��6,��V�.@����7Q*�fI��8���R�ze�ؐ_E�S�ͪ���G�ݥ�\(��A�Dׅ��䝝�\�[ }�YV�߃޹�˚#U�.���|�?���w�k��k?�5��G����W�u��M]D�K��zD`��.���ʟ�_���*�m��]�iS���m��h���+�@$��`�k=��e4���p��'7����"��߄9�R�ސ��E�׿�؅��M��11�rHBEr�ƹW�$U�ة��	����1���	�"m`tWy��'��>#l�ؽ���6>ߊ����j&�E܄�0{�o�Z�<]����+'�"0�����&�5�`\O��.�K
�]~�n�Q`,�c=RP#�Ѻ�@b��}\:�JcXՇg��Xl	��ιߍ'��ʻ�&�8+3"�.a���"�����wio�U� �Ї)��JC�����H@�[�Y�C�h(��JHR�5O�
6�L�6UQ�T��e��꽘�^��F=���:O�W(_�ɻ��2HҪ�k��j��c�\���E��_Y�b�WaE���I����?*vIB1��%+�v�7�EK�v�8Fh(eD�l��t���?���fs������R%j�ߤ=hT6?��Xri^q�1c۰�2=϶�z߄�x�i���aV�c���ON$M��Xg1�v�a���Ç�n���QQ�1Ƌk�O��x8H>�����
Q�%9w��H>W�OޟU��)�P�|�qn;Zϭ1�mt�2�l8�xN"�%���n��
���M{��>x\zV-#��0"�k�нH"^�[<�����������