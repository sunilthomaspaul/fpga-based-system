XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��R�	9���',�,��;l 
�q�R����n����R�}�����f�<�U��da�rv�a(��z*U� �;]q)���.~ü�~�{�l�lf��;x�<C�PI4�=G��b�a1F\�Pg��jQUXj���-����%��#�-T3���n�\�t�B�c���q1�
!"��J�oNߝg2?�u^0j�X $�t��F*A��~��6��	,lt�D������</پ�.o�L�	��l}�#�����m*�<�\j�����;���o�B�����!��U��$V�"r6|��YT4�1Q](��NT��M����K˛S���Ĺ�ܓ~�P_���V��D�]$В��X�4��Ƌ�ܑ�S)�\S�x�u�E�PG��/���5�z<�{8�u�����^��N�τl#U*G9��gA�㼃_Dyl�11E�$=��{![tY����g(�b�?,��^(��`6�sA�E�mf5#�ZK猸��L�T���܆��[NB\3���"MZ8�D(ca��U�����i�l��tNl����Aqϒ�a.ا�j�˶{!�:�D.ߺ��������<����H�C�v��2��z^�=�qa��d�3g�0e�x=е�"C�	:�*��_6ʘ��wYVŃWX�&�-(���"�jI�BG���&U) n��|�`9�J�.��f�<�1��Bqr������K�e��琉/h�EW�3͠�'Ik3��C1��� ��DAX�ϹXlxVHYEB    fa00    2c50���Y�nks@����OI���C��a56M�%�e�eQ�}���VW�nA��sҩeB[�}-�X�:��EG��K|���4�MsVԵ��O��Ny�p����.s<���L�ǲwK�Jz���G�l�\qZFO�h�t���V�܉��Y۴�	F�o�� Ǉ�اE��%;O�&k�	��=���k�0	��0m��_Lq�S�ﻦX���!];�_��g��r�� ;����F�p�(`%�·��dj�e!_�^0ʅ�]��m�}�).�L�/w4��B��ob32]i�PW�io�����G�[U-��D�i~�ӎ�+��%�F��p�
�ѯ�tBHGj>�u��*SF-���&o�SV�'�bSV�-�������dVO3���"A���m����kY�UQV��&�C3Ʀ�"/+X�݈��Y4L�/���E�Z�r!�y��o�ǰ2����9�^ȏ�V-AS���o������[�1�kqm&q��@�D2��.�
@kk�*���Ec���!��D`�;T������r�h����񦃕D9�ps�mS#�)����+�=K%�`>d_V�,��q��*��z����#�����N��H���Z���2��Hl��p��f�{�,�5 {D^�-Jr8խ@㫽��f&KV>U�Q8�j ���x(��e�a���iՀҟ�K���4�3瞕dhO6轊'�8<��)̄��;�M]1��!���a{�Bt0#M�ƒn9��n�#�A�~�D����L�:����Xf�#�l�m�s�I���LҰ'�_ Ö*R�mV3}���w�A�gU�+n�#�R�4�c(���"�)�\nv�B�zV��S��=�0u��Q_��t�Ϗ����	�]���3�Q�f`����C�rIAM$H�)btu�L���/>ۛk��2��aW6��G�ɤ�<�����md).���#�g����K���[��^��1v$�^�"�jZ+�v2��lu���X׻�����C�@jV���
�
79yM�|4(FV�����?��:�&�.)����ٹ�q @X�HҴ�	D5 � y���7���%k�>�U$�gi�#Rxv��b:WG$�yc�a.�ė�(���7��uz��FZ�&g�l=��l!�L�!�u�
y.�l�����t����|�Jo����Y�M����T۳��~��%w�h�ɪ2����@�\}?�o� 	0a���9Z�L���ơ�p;&�.nAA�irR�Rm�_Ġ���[�+�����E�4g���\�\�B��
�׵9}�,���ӥ��Ȫ�?]�!h��h$7�/"�@S|\\�>�����ղ����@mwY �8nFT����vx}����"Ih_����	v�c�f�MC���VpwUA�${�o�T�5��'� F�g���E�oz�w��%;!)�-sO�
2=A?*6����p��~��tF1�~M]�
"�ջ��s�l��΄��6.��"8�����e7�\�P#7�ϓʴ�<���'��D��i����Y#���d�j!%����7�7��!�s�d��5��Jƌ�����tT��M9�^#�s����L�`x���T�S�0;���D�^x���0�8�j6W�� �"7��"�U�P���ke�G{��V��A�AQMߙ6���`1?N��!!�Q;�LϬOŸ���A���ҋ.�Z�$��Oޖ�B�h�f#eIDL\/�ɺ��5�>�O����n��n�� ^� P���v&3>�i�_'���R8�@�&�١v��	t���ܗ��־I�Il!��]���S;��-;�*2g�u<��3�a&v��vڨ	�8�G#�P���D��3�%�:����)�i�J���y���~�K�Z8�(�����L�d.�ޅt6#�%�ѩ��N��Eb��I����_*�������_:�����SYk(�� T_���PfG��l�T�	�U,n��`yD�1GHp�\�%4\���8�B��&��A����e���.e��S�^��j�[oC�	��jV�ol��\=ZoЙł���&����0S i�GI��Etļ�<��7���(i�鎉�*��m�>λXE����7�=��{�'ESm�c^QĚ���̠����<��wD�W�Ҋ�h[z��)�'��G��}1o��+�\i�2��)[��Ǥ��j��$"���U�&`J�=
J���u�ݲP7�W�Q]_i�#`ۭi�8��<9���> �Ŵ0��b���ٽ`ѓ*Y��Q��K�p$�C"�8�@־�����i���  ��w�8�K!������Y1�f��H�-�]�����R1�Z�>V��ZI��z�Zn�k2՝1OF���-� F��x�H��K��rI�����<ɯ�T7��#��H5��\�+��g�돳�ڲ��s��! ��#D����B߉��_%k)�|�v���55���A�ӵr�$�Q}Oih%6T�LvGI�+/��`�@���q���[�.	�<���8uߡ"LM�
C�7�c�$C%L����������@���P��7�c���tM�b�4�J聧�l�PT�����
����]�O������N�bӅ�լ`�n��*�Q�U��څ��Uʙ�N������S7�lNP���fB�����8wβud�A�p����I@�/�k��3��y��R O�ћu�>���o,GN.�9H����,~8�B���}�W�X#�AT��XNO+�D�	;��n`N���Jh�uj�����1,^��%����I�71'h���Y���Krɒ�x�.���Zn5�cb��D-���˴JX��I0�	���j?�g��L?z7�o�@Q�tMo���m�kg)^�]����`@[��-ǳ�ǵ�leId�7�W��V���d����D/�I,�D�*��,?ΐ���8��m�	���d�3�-�80�j���nZ�m#=@������Bc�Ѐ��S��l5U;��b��y�j����O'Xy�{�G� ���Z�~�p����Һ��n\l	N�1 'B��x;?���~<t��������R��
�=]�|����hN2���"���ډ���W��,Q�D@EFt��+����ڿ��S|ΘK<"h����.m0v�Ȫ_GK�����tA)��8�$�{��@��Vկ�*}ݔ�.P_v��'v�O���Vc��$܌]�����P����_�Yٻ��������hg�l-lM�����Ԩ�X�a3�Bxf��6��sr+��8R��Z�>��+V���u�QL	
�1�(<��5ğ +��?���)�� ����eP'�K��9����{�!n���^L�����/7���Yp�	i���%��s����Ƽ�f7��x�YÿwW���V[���lK�� w8*s��
vR�������C��|�����Ҙ�5 Q¨���*Y���D�~%�k�����[N�������9JX;*�t�u"4�-s��.����v�(EJ4f2��\\��j�~�1�Jf�]%T�;�a��1	"c�[��8kت]�8?�����t�=�!?j<=��^W�q"��F��Zuh��<�d������ې���k�yK�~(���i��c�g���?���!�@�3\�U�����09L�{�ə������r$��'���g=*�\o�4�E�@���`m �q檈��H�V�T\��[XϒAY��7���!�+@P�?>h�eCsG6P�|\��8�s����$�69�!m:��m͡�x�Q@�\"�����I�����Y�C�y�k��Y���DL�'f��1=|�ܹ���㣨�f�M���
��n�rB|���C^V���{¥-����	����@���|՘c����h?�u͟Q/m�	mo]��g�.�7��k��p�I��p+x~�z����g��ނ+�.�/��o(8�P	�����R0�+�� �/�32�]AP��@�Q0�ҟ�.�k��
��L=�*���P9&��ɂX���O�!f��j��$`�J䬈O��*�z�Q �'@ٿ6S7������M���%ƺ�˳y/L �7ۦf=78?�-H\���Y0�@H��ТM,�usa�h�lt�9e�T�p�3Q'�ؼ�S~5��먈2dp�Ђ�.�����L}�푲�w�A�fz�Nm�=�pi�=1u���\wb�`w�zQ�o�s���XC�K ���ӟ1����p�����jZ�$J4�xӟ��x��ˠ�88�u�Ri�/��CPq��Q��fD�C������*1s�H���y�� ��o�Bq���3��u��އ�l�O�xMt�էv��g���S�> �'Nq�����\i��!��k0
��=�t֧�I�X����"߯@)�Q�E�e�Q^�}(O�Leؔ�X��1(�;)���	ޯ
���Q6�֪|L�zu�
�勤�#�n�՞�<"�=Y�_��x쒆�n�R
��=vZe���Iu�]���x��,������� 7pǎ\ʁ�X�)"ˀVK�F�	,�7��T����H�C�b��B�,Knk��y�.����U���%U6��Sz֛��UW����;�:�{�D���O�gء*���D��:������}s���$���P�Ծ�ey�/�蓸l���Fǒ�����b����ԣ!g�h��T:��4�
`���HO�ٚ�3��o'$\�v�NW�nV`5���6�|zH1A�[����X�(��ul��X�$W
��X(�܈Ů�FnNK~MS�A_4;1�P�a���֗l�-��U7=�c��< ��!㦰��zdE�S��nm@z��5�	nP)K�U�E�QW�ц�{�6�R���W\
����ms�l,H�<K��^�|�(�y�I��\u$���+�X�c���ػ�9�G��P#Y8פ �w���CS+�v(>�;�m�А�zYV�S׈$`��!x`t�e��ഐ������`=�iШ�����M,�XџJ�}�������w�+���_�0Y�:r8?M����/A+9�vZ���m�{�+1r�zip�r��v�ݫ��tIF�	���+�C�	�\|�Zz�>�by�o�Y[f/u���l�2�����ztn��S.�Jm��
U ?~x�D�x�Bf�trD��DmaY��'�xX��5v���tWW��P�4$��a"����Nʬ����.�;���5^��&Y̿~u�(/"�ÎBq�-���G}�U8����?4o�Q�9>S��"�B�r��P�'�呺�Aʼ(B0`�!5�0���N˨��8��6�uK��;[�%UR����"�)�[Y`�_��-�%�wX�(���J �|��.��?����������
��דX�o[�w��%�l�������Ғn���q~�u���@�:����r��zA/���<G��ȭ4��X؊R�
�|�6��e�]w0��u0Y݊�B�X�>�� �#�+0�2y�y��c�� ��:u�Č5{�BgU���W0�^�󞪀g���k�<q;�z��V�bGH�%*�G�����,~���K|��~� &<��7����Q`�g}^���䑒"O��F��$�?V��b� ~Wjzc�W�d7Y/KP��ւpy!b5m�%TGw��:W���$�I�5�����M����_��t��/�r��%��X̦���R|�]-�AH�0���Xj��L �<��(�����߫�|Y2�����	9A���+�w�5��6峦��ǗqY��}O���>:|��m�?�>����-�|F����g=����ۆ�Y�B"�)j����i��ׇ��ZD�j�Zm Ts�\Q`}VU(-�>O�usv���*�Q×�`=�V� ���+�+��F�(��"	����-ج,A#���n�Y���X?�[�w ��Y�d�ftN J6WV0�G�Jy�bSk	�tž�S��8���Ě�ࢸ9?k��+��9ܽ���K�H2��~6g�,�;⇽[KE8�>KRe8t���Ck��-��@����� �a&� �Ia���D��X4�p�ķ�]s��"e��S����&۷��8��VN�+�X��`.�I��KB��Ҽ3=#C�D|Z���͉��T���ry�d0b��T��@.��1��N�5�ds�����LOO��
I~:G-F�b N�Y����KdϠ����>��������@I�cY����e�VJ�".i(ɯr�杈,���ь�%&b}9Im8�D�U��¾4�(����}z���<�g��-�O�_'ۯ��+��.9�)�i�k�E���ח,��
���Y]�jO׮�|����i�DM��*����0�k7�8��5��(�<�m��|V�.M��������ll�6����%�h���k-�&_�X<48zTa��A��3���0��K���峆��8�]Kx�����I�%�$�}O]A����c��e��6����,��<#������&"m-}b|�(�70���e1�vl����[��l�qW�w�w}[�k~}�t�����x�g�!F����[��j�����
"���	>���[)j�9?����)��g��������]�oj_4�mM�U�;�Ce������v���v`S�� $��e��G�)to$��{�\yN��U!g,Y��6�����́le:nI44��-q־���4Q �0n�K��Mk��6��)_�C�]1��9�B`�:x�[���j�*��IU~��Q���hh�I�����2^� ���_q)@k�9U��bͯ�)�4���lQ�,ſ\��$���3���@HM�&�Nޛ�	�79�~n ���yw�ŋ��醑���}����S�#悽�j�xy��`�4����\���_p4q�]f%*mE<H ��T
ڛ�F�n�![p�l�����F���3c�� O��)U�Q����͏���׏���b����<�E�d�*��G�c\Z�ҶU��bb��"�qة��)�`^�o�)@�g�쎚#�}���О���'}J����2�Ip���ţ���_j8���[�]���`���.Q�A)���1i���j:d�؅ 	����|�[�Wx����>��a�F�kH����X" �a��rvh!�Z��,!�_�Hx�9����	)�g@b=!�U��d�B��9ݰk��^�Ϊ	7-A�^&��� ����i��tWZ{�]'"JA��/:<O�L�f�5%��ϣ#ika����FF�!gY�qip��vm�۰��7��%Ñ���!�T�L�3Z�ՄQJ�!S��5H]�~�H4���$���Q�"�2�D^ު��^�j���C26ƈd~��Z���d���U@�B�0/���x4I�.n��_q�+1���r(�F�ډ�"8������+y�tF��:-y��߸��{�O�>��Fɯ���x��9��Z��X�&����x3ZJe�q�j�{~�?xg[��R�:�U�5���B�����9_
���/�xJ*�TNS!M�����ʛn`a��R���.Ueq�˵��J�Ĭ>�7�g�U�&~`;�Ѩ/t��}kn�d�js�<;����O��4M�?��D�3��xU�D�y��D%)�׮5G�9��vj�v9�1JQD�-/���P�	�J�u��M|s'5��n�~|pE
pl�sA�]Y�i�r��O 2/���t���o��D�i+���>�{�x�P����Wc����4_�̩}[`�t�J��P�.��������Bz��2�%��J����U�Lsn>�ڽ}��N,�e͌���L�Ȓ9��G���+��5���������2`
Wy=&J���UI�O[�˦X�\ OB �t������ �c�i9��G����}�Kt=�ڬҶM|�i��g2O�G�8�n��%��e(���l�M�4��aB�y��m��I�~%�w~Z�����{�o��赈�d��6��5���o��{:G����n����NU1��C�O���"�eO��O����������~�p	�B�7�a��@���XIʤ�φ���j�"!p�Cs�K�PO�o�zrʴ�\Ώ�B:�50���I�g��N4��Sڂ�9NS���2����qb{$ثYX%l+SL�$������Q������{�f�����-7�,`-Q����F�( l�ʳ��3-��[!���
a�١�x-Uȋ9��Kl9��4�2k��pf��e����I�� W�_%��7����LfV�H}^X��45�A+>K. ZdA�k�-f&$n�7F�!��D�c;������r�J��W��5cQ�����^�h,ZMٿ��v�1�"6��ʏ�%�d�����X�%ȩU!R�&&����������m��Y����;�}?y��@�`pe&�dF��Л��<M���;��q����:? 	�d��[kk���oė���8�g�A���X8f��_���h�J�Z�D��-��/Z����
�a�"o_r�D2�c�0d:�Wsν�Z4S ��!��s��P
9qqǣ�Y<��+E��M2���ݯ�ٞ�q�Y+��J�#�j݊�Ph��jB�Vjs�hypU
,+�i@�-Irf�?w{��)&�Y��A���rQWZG�����Egi��3nB�3ȘV
*_#�t.}�Ri�f���hY��.�~eƄ�L�Xm�*i����nq�&��8lX{·'�:�Z/;2Ё�;o���[� �J�QZI+{}�[�o��+�F�^��S�d�=���Z�n����D��%��` ��<
t�1`�[7e�zv^�؄z/W������c ��/yI�����L8� M�>����t���ό�?�K4%ej�ڑ�MH�(f�>~�j�.Nw��-���R'��ףH՞�2��'�D3	G�������*�W����hl�?�)4�?I�;��i������|5�m?VN���@�� ��>HY��;�� a�j�?G���P6���4b:L�	 T�U�[�����:��TO��l�^���U�����[
h̔lx:����Bzz*Z�Y~A���P�)��	_ZG�~iv�B��)TY,���ٮֽ	@�U�>[	3���xVe8�8d��7�3+ץ�Ed�A�wzB8Q@��J�5�L�<F��" �J�^[sc��Ϣ�3���3>��P������pa��0 ��n|d3�ࡩ(�����J��>��A7�Խ+;R{t���@5�`F
�Ħ�.R�[V�\E�����W���#j5��vͻ^*l��n���oD�L��`��.����Y�P���s��ݳ����;ֆ~����g�X�_���9�<g�a�n��f��z�Ms&P]H|J�;*#�L�{k��+���-��&��]����?tq��'�TF��B���w���!*�3P�y�#�
E�a_��f�c��	2�R��!���3�iD+�Q�}�k���e�YN��0& ������wi �'bj|���<�.ffC�����W�6�8��zmA����;+��  �dq�����,�*���'�&D��5T <�D=���>T���ś��E�"�FJ1��*�7\����{�l��V�?7`Ü��ew�bS-���䅇}�wB� H�a��}�����Ym�,��	��H��s���px���T��* ��S�k��7OC؜�zTqi�g�}B�_~�=�M2 ���#DJRI�����Ό�7;��w��4�hp;s�A��9�C���k#ݻ>ɪ����)�M�e��Ɩ��B��4]Ii�\*2S�u*8������Z|@c�7V;k������c��@���4e5��@_�3�L����E�{�2���o܃e��U�s��4�NR�����/z?����88��bRe�������8�v�B7����鎞�7�u�>$�t��vw1T5*�t�ߌ/�'��Xx��Ċ�����Ȧc!��J1?Q�k��y�����1�o�9H�4]$�
.��pcu�bY:�i�=�斎��R��� f/�a�d\�M����xM�dG���	q�Uȍ��0�!��Q�i:�a.al��'A4�������&�A����H��`N��ߋ�
:K��H�1 ����殚�e �d��z�m�{��[N�h��Cr�Y��LEX>�+V��� d�g"�6���[�l��',�� "�V��w�r����z3�9������"��6Cpr��!�*��%��E���Z�*7��h���>��J���Bh$��}�O8��_K�~��^��(��ᤏ�Fd�;%�8K��A��{���b��a>Ξ�p�P��2"a���ԡ�7Rd�fۢ�J���̳h;�R��<��I���!��<�4?�;���^R:�rkj!��8�UX���~.�u(���ܼo�V|�l�h�'h!"Ɇ�-cu����*����?ɑA1�����2mk5W�q|VHc(U� z~��.�p�.���k	�E٩�1�>A�S��')�ݦ�H:F�S�Ǧ���)q3�B/�Ԅq�0y�+eAʴ�?4�xϻV]�.㗔Q��{�-���~�E|s �|�[����R���)�8oA�>���d�c�='Sո�y_��%��׉x�����ש�^b�q1�7R�Yo�0�I��У�A�⯦)A���䉞Y1�W�4�$�C=���q�dę͵�P�2ET��v%�Ng�pbI���H�[�H0�?��L���.1�{�1*ш�X~.���<��C��7�h���p͌,�*������v����X�6��#Ѽs���6�[l����b��P����ĵSj�~����(D�����etmB�(�������I!�XG�4�*&���w���Ĝs\j&ё֏M^�9��Yu�>��ӭ��Q\t�sM�vԢj]^mp�~"�[ v|`J(�ÝecU� �����Sc��ߐ��v���y����i�XPV1��?%�$�|�v*%�hs��}̨�}�񝁸<W9]��>�Ł�,
g>��Z�w�m����m4���!��]�"����q�h�o����?� +h���]A
�X!�}YF���32���˥�����j`�#�U���Ӆ�<��$���f ��W&���'� ���=!^�낖�I���Иi�7YS�XlxVHYEB    c397    2030a5>�1�Y�{B/�D@](Q[��(��ov���jZ]�k��Cmν�2(���y���i"O3�~��O��g��	����2&Q�ȂB"p�ZE��Z4�_+�;$�yi[��&���,�𳌹��?�!(�=h���v���e�Y��J���Ն��m���J���YԬ�R�M9����(�Z�]�()*��0���&4�U1����[}�(����O�X4��;l ��B�
 ����S���Cє�Q.�\N��u�0b䞲	�-�XC%�($\��O/��3��O����Dxk� ��X,Խ�6�b�:��N��+�#zʕ��m`�<���#Hƺd�!����QbWQ�˄��H���dE��Ӷ' W8���0Z�+"5�Zb�����61\?�?M��LLV�V/gP*D>'��VBw`�+��j rB��
B�Pz�8Q=�7�-�&_��z?�A>�;33_��RG�L/K̴�� ��R��7@��r�_���6��W*`�`�sp�gG���RW'��ߧyW��ˀ������͌`5h�#'4����,�w5�g|���*oS0��V.�q�>@YH���o�/��[��Ol�X����%�^������=8���O<ȅ����e�uƒ΂�o{�+�����~��L���2�͔6#�d�'[�/'^b�����|ж����L�$�:l��>�ZP0X��-tIhL:3��R�����jvv��N������D=�.��Č��;�Q��L\oZќ2ʹ���g��2��frv�0"�z=ln�|���F�xh�F���Q�j��8)�N���?����"(�%;:�d�$��O��9��[��b��~X:�'"an�z!}T�͋QOA;�0L���*\�?�\�+%�|z�;�n�.���ϬӤщ/�7F��k��og�T���Cz��~���Xp4gj���:$�U��� ��\��K�sRF���XP�^f�?�S�WO�Fy�3�G}�b���+�,��.C�@��u��þ7�uH�����᱊��MX��	&����s8N05������RI�Α�����	�S�T�ac
*����T���{� !R��N�\a/�:��JI��B@,QG`���ϲS��͕BW�����QW��]�P��aQ5�5��]�^ŉ���mfJÚ1n���L[��5����j��<#� 7}�D����n 	T�;ݸ>@�okП�k9nl�^shW�� �IB:+9���j��AG9��!&b��h�r�G���*�X�ʿn��R#=}reG'l���b^׽m񂲳���C7�)�u�P(�� xt���M��c]����O�V`�MJ[��狇n!��$��*��D?�
���Բ�������:���s6��Y z"j7�/@e�S���rL!�� NN���A|8 ъY0���b(�)d*��j袺�A ����xP�ׇ��.��"B� �X��d*3��*��ƶk���{��51���q���C���������0��R�og�߹�#��m ��
U�P�u�>���/Ⲇ�ŇW�LR��@XK쩡;Ѵ�+i��d�j�AK7�C ??uA�/����[�&���nA¶����5�N_����c�*���k!�fG�����Dj�|�������}��{H�"I�~��dA V�&5x�h�����Y�C����H�h�+aYO-��k�G ��('��~a��p�ԫҐG���`0���bkh��á��YC��zc�4��Z@�Q�`��QC��oN0p�9��|��(���jQ3u	��ý�A�<�zt�V�u��r7�~�3�ʎ1'2�ؙ�	þ����~Z��1����C≘�vA�0٥�|�E�m��F����fR�I�v6Qs`i{�nʼ�gM0e��y߱KG#8l	��`)�
t�hZ,HRa�T)X	��ǆ��ŷS@7=���dA�w{Q�U�l*�!T�I5����w~r� &�Ǔ�N�¤r�nD�E�/�R����x��/�p���-��w���Vʒ�ʚt%�e�1ʋ�0��?�5^-h<,
���5�׾�>\��lfۊ��\���)�E��n̞rg]�P�ۿK�)���������	�?!նk��Z�܉yo2�;9����8�|��Ԁf�mU��q���ʪ��#�@�aL{��H��	����F�Ni�M�wU�]/G\��\Wɤ�V�^1ޕ��|�u[�Q`��v���}�����HA��{s}�5���I��z��{��__��䩽E}<��*����՜Q�O�s^��B��J���j��#2@�Z�LV0��O=!W@�׽QO�R�an������(�eg]U�śRXS+����Oz:R���%'���A൷����)�!V����vl^������iM��JUV��&6�YOs�)v�b���P,T���A`��"G�����՘x*�} ���Zv�j�Y�e�X�N1U��D� ���C�*#��}@��2tU��JO�C�1� ���0��jO[��޹m�`
�2+Ϟt�ǔ9�[EyVڱӲ�+c�Ωk��CB�_��o%{�Pm�C��'�G2囹�ԬB(�<CQv��0�-����&$�ϊ���t�!�ڋh���EP}}�r_޶��I��p�{ Z�8��m<KM��e=��������jI�8e��<�:�OzYg���-��PHfU���瓋�����⥀����c<��`?J�4iю�R���2{�o�)�2�,�+�2���xm�fu��/&��{tO4&PhF�F,t#0 ��/��e�	-�+�D(E_T�i�ם��=�y��E�!k`oӾ���V8�L��x�s���F�{�#��Hv��Pl���_�����I�S_��lBW}W��1tWEu��!M�4�����H�3�!��PzI ����G��N�S+Z����� �~��FA��I���uΠ��/�SQ�M�J�����������D�C���8��DXJ0�dĲ��O�MaިV4ז��i�HEt���.t�'�@�V��:2���b�������f�h�X~��U/B�%�\%�w�z�aJV��65��v��S��
f~+=�6����Dġ��V�z5ӣV�ô�U[�zH/�0�1�yh��Q���J�]~n��C6����f�p-Á�Ęq�k�t������W��ʀ�%#8lfޟ����y���:�NC��k���-k����"����E�B���$d�{'G՗��	�潜�f����fB�h�.�#�Cj*M��+s-!l3��{TT��<2�q���ۈ��MN֖��
��}̞�=�c?da)��
��H�Ʃ�O��7��l�l���y$������������?$��\�JL���Q��u5�~�U.�ٳ턾�g&(DG9��M���i%��ά:˷���
�ki�K�%�����-�$���laCM`�-�rԥq��!�/ڎ���dI�P\�#�ecTr$��V	��H��51��q�:�Ӆ��Dg2�����~�.�E!�P4��A���8�k���Nk���h|��������O�`\�����F-�Ǹ�> v��P	��V���N���ʥI��L���6hU�)����g`��3�cm�*���������Ä���8e��fΒ(@,d-�V}ec����ٞ�P�m�Ȋjkq�(�s�i�ר$rCGӗ͹H�-���%��'���[�J:�oĚe�q@9o|����̅G��Ff�V�m<ཱུP�שRr&������ٌ�Ё���0/�ҿ�W��N�JQ�~�|,��?�|���pq��@�þ��R�LL�%>�� D�T0>@[�2�kO�~/}J��E}���o��4Tc���2��|�����u��2�&��ltdc^��Za$A���bd��毹�c`��*��_�j'�>d����������1�<���J&� N0�g�o.@�Ϧ2X�6���)����U�8�P7�fA���٨�P�B%'a ���>�GXd��^���v��<����a�����_��\]{�C��<bp3���7�.�v��g`�FÝ��\�� Yߢ�-Y�?e�dJ
&�J���]0?bC�0�%��N��#�a�Wj1W�M�9n�?�'����C<� ۤ��͟S���$�j��#u���=@u�z�b3�$Tm%Lj׹��t��~ѡ��7�!v<tr��~�U�?�*R����V�KQ��	�U���r�a����.gX�%9��Oʚ�J�Ch��dj8��vGmeqn���!���V����n����o��5+�p�0A���C���r���9����MO:���4!u)��c��Y	��l4G<+x��L$�� Oy�^���N��_
 r[��{��Y���6�u���\h�yq�/��������7��IOa��ד<��Jm3�8�S�<����Ҳ��s�����-��P���PڊR,!����e�e���o�'�����R�7��h�u�V|�U��(V��B�T�o��~����F"��RWyF�z��v[!Q�M�E�)��N�}d��ԯX� �[�t���݃���L5��R�$IK�fa�)�N���xvw_)��҂P�f�'&)����D�'ږFˆ-�G��1�ϵK�|�l^rru��t`�e0��0@�B���yÖ��(U�
�J�	��Pі��ϟݪB��t�;Kxێ��2�\���VlX�)>�����^��rE���!�bJ��$y��R�>�[�*W��tݑ8f&���Ǖo��{��6Y�������8�4��t��aq�EC��ۛ�R�]R��Ra#jy���E�(��LGR���;��óћ�QZ�L�Ϳ���B~T�k@��0H������4����:�J"^�<��S���oW�##w[0@�=y��ߧ�X�{��몫B��!�P���Yx?�����x�&�M`"x��F{_�E�AfC���y<���F�����o��^��x��z;6��9��-�9Kv�W�?�eg�eȽ�du����-�rP(�X��W��I��%S��� ���*_q�_������V(����áz�3��V7��ClA���'l�f�w���p(�}�`��a�	���]��@�| bл�(�Pi�"�$'��@��,K8m�Ec�_�#�Ϋ��K{�xwێ�d>�L���s����E�
�ǌ ��ʜ��tv�C����F
�v��p���E3p��G��j�v�"��<���aI% `��!�x��0��3"«���S����G����'��W���s�'=c�<��C�\RN%h.A	dV!�$���OC7�k�����eM��k�犿�{�C�@03��@��ȚۅdHĞK	Mǖyvw�@��'�-���P�kO�h�]�3�{��wL6y��0$bƌw�=��k�����:X�o޽98Y�����!��~��T�_���G�8��]��۝�a5��t�%����j��xc��۸U��=��9��U�'��|"��]p�}F�1�NN�j�&����0U�@�v�i��p�Y�꼙�tF}����ƘS+[�h_ܓZc�/�S�P��A�1�����?H��G��9ՠF
W:���_8{�Ї����O�����y��
U��)��hJQ쨌�%l.Jn���jYJ� ���a�v�0ǂ�%4&���Z1��dp���dR�H��y����<�oq漮��a~��1��F,?�]�#�ͷ�	aʍ�R&!K�T��R{�Oj�,��[I��~���"�°���B�վ��8�͑,x�
:�P<_Ǟ�5����V��C��;��zZ5�����F�|ZP}��_����Iw���	�	J	ʘY���M�cџf[
�=Jd���D�o�.v�}�U� �����I�]k���\r�5���9w� �����7^2�Vˠ@b!I'�ۍ��@t�Aa�R5�y�`X�or�pgX -/����?M_n��c��ኲ�!��9��y�cL1F&��S�@[<�4@�I����8�U�E�W��X;�R1Ni2�h�X��ݷ=A�+R��������|��e��Ep��5�5��{:i�1Q�V"��|�A���Zߌ:��eG�B4��[�`���A<H%����ܺ�Kv(���y?�Psc�c�#�#E��
Fs�,��z��^% �nZ�w�����NW�����y��0i��7��n�S�n�y�L�n��eQvȿP����cV$`(�Y�U"#�X�BݑW����~U����*�)Q���D��bY���N�R���˃䫗�J�����j�V����b|���4(�sCҼ��8�X��z}��bz���O�-1����� �NN`#1;�Z�X�Q�sZl�y���a�da�C�\�9ѥ�y�3L�{��:�7vS�!�IEz�NX&bR�Ǟ�v�fqB��h)��G�F����.��\��u�\��#�˥�_"�����훡OA�"҆��B�P��=I_�aY��,l�0�_=�C�Ĭl����7�C�wBJ�9�[E.!&{�ѣ�\� _$��8�y��hY��u?�� �@�2Û�s�p;�k�,h���
Χۚ�g�ϭ�վ�Y�̊55�?�&z6�ȿhj��]�Eu]2.o3�Z/�m*��b��m˯�C[�[� dcM���w��T��
9�Fm"%q��(ѧ�
%��f��O��U�@<.2X;Ѱ!I��2��Ҍ�ND����>��X� //H�9����0��˓�5�����P?��#�Vc��9�K�Ћ+VA����d���ES��VA�;�L�t��)�n�����k�l��k�,��<����k���7+���b�Ț;o��u�6�nBk���\�jbY��P�e��tOY\*��@�M򵓊���.:�Ugg�$���X���M0鬍�_�w� ��pq�s3o���������ї|X�9�h:Y#�zn��Z2;��sճƬy/��7��e�菡��[	��Ӎ;3/�s�HN�P��^K�W��<���l��bQ/��H���u^V(�s��fwy�#�.�Z���|Gr���V�r��i|.R�Rtݱb�+F��h�M�>�taQof؎���6��)WF��g�N��tM��W&���a_.W���0�C�~��pK��[�^�_.ǚMcoO�P�� ��� ¶kf�G�̴C�KF��bl�0�uV_e�f��CЈQ�F)���7�Y��=�[�����־j��2тO�=�ӯ��6▰�%�a�zz��5{�w��\��!F>&LY�3_M��3b�|:�������V�Hu�a0�cJ���B�t'�1%��ضߗ�D	h�aJ�F^C^��j��]=&U�p�O��z�U�)��<,`�FM���0)�t }��Jfhyg[�W�h�Vn�0$y�@���dkd�|Ӊ�2�z˛m�֚���b�f�%%���5L���%�hI����.d4;4�z�Y�%U����e\��)������&}�\��Ke&l{
�$}"���	�ѡ�SG5ZG��.��
���Q������*F�����'�@t�yy��Һ����������Wk�X�#�DMgY���JI���~�*YQ<�1�� �NM���@;QM�/�y�mo.�#��-���w�3�I!b���?@�!_��{L�=6���o}�:#�����S����s�H�}����t��?�/��1�g�L�BUo���u���Œ��ߨ-�U���%�*�,A/ �D�l�@��]i��=`����SC�V8b�*^�ެ�샓A}�F0w�	�wn��OǕpꮍ��Aia׋����d�ZW]4ӿ�FB� ���sA�vE5��F.vl�ήl7>���eE���O*M$��ܛ\՘��P*U�Ń&{�F*��o����m_d�#��Y�pU+TEH#�e`�����h^T�H��/�ԏު W���;�Zw�n�d����Y^��:���b8d�� =J���:Ӥ��ݱ�%���d��;mG9��36K�<;�V����Ӕϴ��JL"l�Jtj��6	��V�&wm�	&4��?����HR|ytH����Fzÿ��6�-o��{�za�n{������h���
�ze�}�3�a$���.���9+��P