XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���_��qom��U��Jh)���J�V-�?K�-}֝qd��<��]GL��/�Ξ�T�:sgIS�n��*5K��=ļ����F�#�<i�_�ݦ��.�4�0(�ln���<��-[��_|��-E�)<=���gf���"w�V�qa��gש�������E��8շSDm����-q��@v�����#�ZV��ɮT `��R�	�\��
����Hp`%�]!����Y�7A2֎��Y��%�7�L�~��B����A2w,��D���,W���3��wl���#��/�Ij�������|PFLo�=���d7��W '�uTƧq��	���r�1��J��|�M%�v�8i5��I���	ς��ֹTa�לBMϩ.����-��80?&��\q$��ՁkM
��_;��M¯˙HȻUL+X�v%6�d���
�ȿ�4�7����"��s�A�U�N-��dCͭ����g �~�sx���Dg�<�a塴ak�:d���2���A T4�A(�9�d��������3����#����.K;��/�4Je�V��������p��p�� �uK�(��)^5�C���L��N��z�A{���9��:��[j>����Z_]����M%�~����t�0L��7>4�8՛�`�<�e�<?��J���������C�B��O��>�x�J�-M�?�|�����s�7���g�+���O��Nu��j���8̗�D֏�e;!f���`U��`���2{C]�XlxVHYEB    2442     ab0a�:���
|�,�4#4��	k�G����@W��7V��� _�n r��D���M�����
�W����Gm�+�Vqr�@�eh��mEc�	 �f ���\��I:UU�īl�o*l��s�=�s&Ϟۿ9ur/�*��F��@b�������ad'��,��&�s�?)�����7N릆f�=r�@���SYy(&/�'�z~����pw�79��-ʇ�P�H���e�4�Z��Vs���>�:�n��T����E����U�XE�f��\yr_E�|:.xWDn9!�!�����|���W>� �A�1"����%��I�Y,0MG�HN�|�����B��c<�O`�3�3�TY��8W��M/+�|��#�E�8����y�=� ����8�3�ްY�"-�|�W�S�F�Z�Q�_�j�M����i�F�"�Я���k���O�I}*}O��A=j��3X�6c�]�~;��p���T�,��.�O4�R(���/ۊ�sqW�fyUZ���|=�/��n%���ڡHq#U�/y/R]�����3���B��������jquҢ�x;�?�z��^;��E�\>+�ݮ�����`�~�UXa���AfAW)� j8���d�E%FY��v����:��f�O�^�j��Xq;�����ntM��Ul�5JM��Z�dRq���
�\���?��!Q�)���=��~�;�Jh�OK��&��&O��i�s�3�fLF�������2KMG�Э� ��bқ��.�a|--��1���-n1B�����/���<��*H�yg)�H�[�]���.�:\�	A�Kc�~]��e6o1��7Uи���>���8w!C�{��O�����#HcŶ�gZ�]����\��(�R_��F HN�TI�޺�8��j6x	�k�W�������@��u<7���+��ucO_N ���u�\t%�a�9.F�t3]j�niZ�a�f����Azh�
�
�}�`u�C4~c�d������c�ݒIXN����ʹͱ-T�$��=M�s}G~�M��*DP1��<���8��dͬD�3b
G��O�R����S���뿤@�j��$��wǳ��g0i�ϗ�g�s�[��ٰ�i��O�F=�9Ր׹'q��w�[b6���S�T�ʖ������������9��2�{�]j�
Xkn+��0�M;�~�]���/6�Ca���8�^���X�ਲ਼6'�8���d(�#�(�	٩PC6,���B+�+.��&k]�~��<�m'�i�_��@�/�����c3vĕM�������)�Ͳ��=�<Y+x�r�]M��g���<Oe�oP)pG�0m+{�_n�磄�d�SOi�g��	z�+n�c�QŃ�L�ߪ�HMvy� �!Fя��z��S$O`E��I��ü�
#����+��<�0y$�7D3h����5��C�*��B�̧�)��m0�%�����i�R0��(�K��{�jhb����}�3�b��������u�m����Go����u��>s��W%����r���6��eJY������B���FU�jަ4�+;i�4�O���|�-B�c��Ӱ��K#�T�>U�yo����� ��b���s ^�̙���� z~�1~u�Ģ����w��f��Mpϟ:Zhڲ���!PƺscjS잊�q�L������|�.�8� �<���Z47�7�Eh�97o��nr���>�}ct���a6H���'wH�����+�[zEy�Q��lȢƭBu��-'�@��Jo�ZTV�C<�\��� ��u�L�!Pk���k�s[��w���Cp����M��E?
�=pX��hB�?2y*�IM@��li��8��ih�I�7E3:>u�^�&�-�8a��2vx��`�Q���� C�^�M���$�V>.�ώ���n��j4��:�6�3�%f^>m�m]T��Y?�Ϻd��u��E�=w��YY5�˼���� ����.z�7{ҙA�sW z�X�W p7L6ا��b��}줙L�v`2G*���sE�sY�G=�6-�}d8�:�A��ރ��c�v�G~Z��ĭ��ɝx8�x�\�VE�-@׽fu��l�IW����fP>��h�2ˑ=B�7M��G�t�Dz�_9���.x�)�m:�����k��:��t���`RFZ1
�ˎ%��Z�]u������^n5B/���?;>�69�{k.�֊|@;pҫ�D⾅��FeDO�u�{#��R��9�D����'��E�[��n�����f�c[7���OQ�q̕K���F���Y�FR+�<ol�^�Np�~o��IԨ�>g')���%mF=��ֽ�`e�d�Z'���S?�N�� "΃"����I�FC^&c2$�!�q��j�_��^�6s"��W̎RkFj3���U��� Ir(ogj����z�=?%��O�y��Ox�1��Rc����@YI�Գ/��u�����s�m�n�Q
.ԉ������7&[��֬�(�~�k�U�� ͙P8!��BW��:�^�s�("[NηAk��7�%��h1��O��HvPP�-�~�ٺ7��J��(�n��O+j܅*�km�+��g���L��z�J�-*;��~�?_�6��!��x�ۮ��j�>��,�H}�\L�&�j'P}���?KޯÅ�Q ��q���I���^r�5� B�\l��+���J�����/���