XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��3��x��\���@����Q�z�|��ӯ���g54����X�X .����B�Ka{Y��&����j��##�m�+�˛Hz�瓙����`�I���r�6�;s����p�Fz7����G�����r�
�Q��V�_���C�Sh&�;^Ysq�o�a�f�L������$F��Mv箤��w��m��к�:���s_�)���8M�&�t.�%iZ}>���¡��<��阣��cI*��Cw|7��@����P�ম"Ώ;Y�ѣ�;���"�����0!�N��1��3����V��֤r`�2Q,7O��ee�_L�G���%�1��r��I�����wȲ�|1���¡4PѲ��Υ��s�:�G:�L����Li��f+��$�6��$s�g�]�ʳ"��)�p�4�����H��G8崰2MU� C���v�qtG꺗��в%q'�;89�.vL�+�/�Ǘ�����O��$/]��@z��j�Q��R�8�CU���LǇD�,>W�8`��w���. D����f��c�^�W`L8ݪ��6���doz	����
܌�g���͈�@���Cҥ[<(���:|
�Κ��}��4��u�[;���?�׿n�'�=�$�/�>��+��T�x�1�{&�U����j9z��-��<C_��xd�s�-��fg+m[�w�d����c�\�0�)��+i�خx�u��B:����<&t��#洚�w ]���i'.g{�6��scXlxVHYEB    523b    1130�-��
����b8���`��yQ�((1��k�R�z��]����D[�Z�97�-T����I���&���^�CBC�n�Y��9�P���E��3�h���j��	A��R	�r�̟aW_/����J�˳�;@y(M�fg���:'�w3�=w,��*�^7K��_zN�����b���DٍǇ���R=$��0K��g�x�Z���xt�Q��Z��*����ǜ�͆�k�?�������UԷ�o7�'��Re��5��Q�#��<�ê�(�����}�!\��ڻ!� M���*�� �jd��|�����=�S{�����?z����ߪ�s
u��'��n��|����3��~� c�D��Qae7>8\��9I����%-B�-�p���w���Ua���sۡ.+F	є�2����R&z��a��r̙�ƥ��X3}s�);j������}����*�9����ԡ���Y�,MW��d�-��/��u��~����o�kJ�5���a�{�0\��O�@���~�*m�v_���Q�*_V��B]���tp�|B�5o�������ح�1>�0ڵ^B|D�D3��6pT����ҕ��+��ƚ��������0�sP�
c�,U���	>�?���dw��n�1tcu2� v��6�t�8���8��Cq��?_QFp�Q�cQ�>�_����=�<Ju&mt�,�[�5k���i/I�D ��D��E�:��X?�ֹl�ୄrP2{/�q�f"���:6.i�ѥ�������Vң�e:
����f��������~�	Z Lhړ��h�=�I�'�P�Yg))	�m�����jQ�����N����@�B5}�zD}ξT����
��	��Q�+�u�1$#]�\\mA����d��.j�X,����\51���c�n�0`඾��D�$b�p�c�</bS�]ll�pkc�	7u����t��l�Yz��� WEmKN��)�c&_
_�=x��Lnׁ�aONh�3���1J��ej���O�o��`�>)�6"�O��3��3y�Do[�-s����������%l��l�l�G�rW����\��x�A���J�JޫX*�F��3��d	0��gu a��rf@�wmj�B*[rт�v9�N#}���e1ހ8d�x�"K0y���r$N����u h��h���2�7H�S�*<�D��iP�"���;|�˭�M���ЂjM䁰A�-F8ptC�uN��syE��W���w�lbz�3��'F������1�Q>V�d��qE�)@q�$dX��.�uF�^���x��-0n�A�Q&!*�<�.#i]Tz�08bl �:��r�3��'�z���å���E�i�#���O�(��^����$���wY+6�]��"Xq�{2)��?�kt��G���ziO�?e���8�y&fi�eݖ�H�i�{lv���z��P�?��a+�$��4�	zO���H�eo���b����sx��J�
��U���Uh�n���בU��R:���������ߣ�:k��[l�&i�@�ő(�@`�0;�B�/	�I�O;Lۛż��K��<������4�@�xC��?�X���v�U>R^�����ۊ�Q`7�S�E�x���4�ye�I��J�0��R�'��@�&��t�7��;p;����bG��9��7'��:���<9͎�,���.N�v�˅��B�YZ_���b|Nes��߸��Y�e{bBi�?��B��־;k ���G=(F��D�&�W��E�КC��u塪�f��}ڞ��NZ�	`��;l�o�o���Ĩ��\�d	`{�����7��0�3����td���4!q�a��)����#��P[�\��;O�gt���}%,_芫�ǜ@� �ך5������r�q��NQ��Tn�vn>�p�����^ӑJ^�3k���*�ȹJ3��L�QnU��������ԫ����ۜk����S��ی}M)嚗i�_�dd���K��w`J��HB�h�� fR��usȱC�U#e��fMyep�z�^���C�A�,,�CDJ��(̊#��n?D \{�=`n�)K���N��T�����7�H�I��W�ׯ`�����-����Qػ�		-V�l�kE����=+�;p�&�'e��:�{u��h�֐x����O��[���J(�sQѯ>d�A��}P��@���>�R^��p6��������'�g�!���"�Z�6
|"��9@�M�{�/�k��ʋ[(��$z��j�͑�}�m�窋}�Wᡙ�;؍e��^������Ŭ�v�2�樏�?eC�����4��*�Ο��g!�̣�~iA�����9,��6o��(a�!2X���ˈ}�`���`F��&�Ù��@I��v��Tr&|�V}��{�`$'��a�/w���J{�؇�|͙ѯ8�L�4E�^����D�&>�ZJ;���(�5)8g�MW��pט���G>���y�<��0������z�m�GG���|��%���d��� ��%6�g�n���8!�� <W�t��������,#�@w�"�nt��r��Y	��,�bL�L�SH�E'�W�rT<�Yn�m�X���&9xA<�����Yܻ��7Tt�,9	�{	ĦU�{�-r�+~a��$vR|�=�p��7ꁼD1��w�]��'�u��	��W�M�+U��۩��I����Y��ǒ��wX"�di�P	TҐ�@A���9�C�n�p^�s�j=:��� N���{�x�oU�l��u^<,e)�x�zsK�����I)�����XA	�?[6_0/j5K�]�$�A�$"�П�l/J�'q���x���> z�2)��҅��cQ�i�e������BYm�xW�>��N�z�F�lN��4KWH��m�ʈ�ۊ`*��'K�	���_������w��2Y;�RA��$c��
p��T����:�������=�K��TlHP6i�/�_����p�#���I5Ro��.A �����Zٔ�ęX�폼VL6[a1X��rS�S�p����&ѓST�>��F0cc��*!id�+�l�O2��NN�{�EKBtbͬHY�r�vh����� �a9���l�$/�B-���c'E�Ud��y������G��Ŝ 
ý����w�̐2D�f�[�xw�l�Y�H�/�aP��B䘩����9�����:�YDQ�o>����r�~*���ܴ
K^>qd5�e�5�E*���Vc��������T�/v${aV�)Y=w��Ю	�4��W8��*G�Z�q�d|-�ߥ��P������%��_�KuL�9���v�A
�>\KQWr2�T��OmVo�J�0��HJT�VP��S�w�%�x�LF�������l�V�Ix!����3r \᪺��!�et���z�d,[=��I1`�[���8'��rZܡ��{�h��S��C<cjݿGc^����&�}?eȗ����d<n�����v(6�msƀ�,��xi���ɂ7�M�i���t�(r�iSʭ�"Gh���m�_���j���$Ұ}��œ��!�e��F�c<Mcs5b(2�2�$���U���]�0y'6� ��~����d��m�D.����pU5�Cn�Ea�9-:u�H$��8����N\��,�&i;�;E�Z��v��F:�H�~#�mo��c�cr��Y��4��su������mG �l >��T � }�m��|z��N� ��5���f��p�8*�$z�7��yEeTߘn*��l'��3�h�9psxv��\io���r�}��ϫ����gRՁz�q� �?��5]�K1�"�����s���<��i��JP�J�5��ZpX�"5XX~��:}��W�D9G~��l�����c�_����S�	"dxɐYPR*aU����6���;�E�Y��*aU3�i�[J�t���x��@!��w�X�'q�%��a�n�ۧ0X���i�6�'7
B�Y}HC"���"��l���D�5����b�]uE�&�L�;I��f���L��tv$���n�L��sh &�0S[�,6�nyU�9�wG���On�4{�M?��+�z���%�3�&����(I�/���l�[�~Ht�� h��n��Ǽ#"t��Z�g;�$��:%�>���o���uh[�(�?�3 ?���+ɂ#m���q�>Ddr��P���#.Y�S�z����ш����N��n[��k�� �&�Şz§�����.F8��!S'��l�vz���4�e�ڴư6I�B�����2)ءդW�ƪc���j�,,