XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���^�K2��>��Ľ�>�F/�2+�h�<~����������{��b�BX���׋�.�s���n�&����ey
��`�"$Z��^�m�V�C�i�O	���׈�tY{�z<��Q�>���� �c�Lab�{��]�3A�85�k�_��ibF`5�a��-��6�y�S��ʝ�� r�I��|U����_� Q W!X�ڏ�xt�@��^�߮�]�/^$��A��~�{�����.ഌ������njH��yK��t�e��] S��ٶT����e��U${�rp�����ꌛ3�_@s���-]�F�fv,�_��R��=zW�?"�5��n��[&+��q��!�
�i��l�?�týTC�;p#��
0�ծ�Uj�+`ܳ.��T�[��A2�e�|�L���Kʩ����b�$�������PD�\�����Y��#v<d|6-�h�ڠ��g^g��"_�-���IMD��U�
���
�S�:�T�����6#	P
S��^jp����@��̦�T_b}�Q30�YZ��Q8o�[c]�1Ӹ<��O(r��	�����,O O����{D�@KŜ�"u�[�]TVh??��3H��╖ k�`�rY|� 7�]�ɑJ�egh������S�Q���:��C��#u��x��]��y?6�% Xĩ~�*jGյ���ۥQEK2VN�͢�1&��R�a��n��啿�;��e�.Z��Y�*G���J;��EL�nT~J�)t������nt�o�n +?;XlxVHYEB    1d01     a201�x�D��x�`ka�R~C-*d��G�L+c�_C�]����{�FW�(�w�ѼO
A7��+�fB*|��ш�;������8³�`��c����2���?4zL����k�ǆ8�Lͣ/yiA����ռl������ 2�?�X����@�-vj����:��x�~:9<G�`��WV��lS�V��' �hB��֤��`T����l2�^dH�����QԂŏ8lk���#��
��W��㡴���t��e�5�M��k=���w0|�dq��	B��֯����E�8����B;%�lL0��9~Z2�ߢ�|��h����*�9�-.�\	c�s&f�j@�����@><��k~�Q��Q�XwVcx�,��(��p��C�Ha�o�&���	�������YL
nCj������ܜ�z4\�m_y��!&%��˧�|�����i���8�m�'�7,���~�X��k�Q������(�刜�贚y�t��KB�$��{"�r)��"�\�F�-#r�j�3���p&�/m��x��F��-��<x�R�
#�\,6!����"�։�'=��z���Y\Q�џ�)���N,��Ѫc��G�㍊(�`p�4�L���w�\����o�r5G��h^�2����g|
�����g�����{�G@��We%�5�D2�I��C9,�I�٪{���5���2xi��Zx֟(�I��$�נ!ߦ�L�[���'lQK�����hy8�.�Ej�b��7�>j�9��=\�:G!3�&q�
��2��i�����^��J��'{�e�^�^f�o�Ձ�a!6����)��'��&Һ�S���tD��D�4���$�a>K������h:�vl�#�'[��5����Ff֒5��/��ܸh���c�;Lhd|$�lӮ|*���Bk�kf�n�p�z��B��M�qO��cY��w�`}�y��Ѽ�`ƅ�h��.6�G�9�>d2�yJ'-2`QUFS�VϮ��j�y���XO)mu���.i����uz�.�2}����X����V_`��-(j���<.�?�(e���ϗ�B�/��Y.ro̓�@L��z���დr%��e��T�I�%�����t�7���!�~�Z��M���>������������W�t|ְ�� OD�~����^� P��.2X��xVI0W�4�T�J[�Ƥ��|���k����_L�_,Pܐ5�B.�D��nP�t��(8����`�4�w�
8��W�Hq��x1�U�f�U����x(i���¥�%�հ�V����#!j�u��]��(�ܿP�2��~���Y�f���A�c��]��K�>�s�����{U�L2�������K���qǭ�,�ZgϜ���ۢDu�ŷK+W!�L�]k���;�KVJcJ�1�'��?�n�+{����Ȧ�ؑ����?��� �o>{YG�(�fv> �J?��-Ϸ`D�H
�����
[�K�3�'/�%��WW����$�Ŏ����x֭7��״g;sS�rP�z���}>W~s����=
���m�Q��	�p ׀��'���\�P�F��ԫ5.~�J:�)����&��b�,�l�����*0$���/����q��j��47^V62� �K����� �"��Ui�����Ƅ;N�"�ьs��(+��H��)��L����feמ�m2�3F��6`�����g�h�P~��rrM6��!Ї�@T���9LA�Ν��77o R'
?�J1��V���� �� �.�j��;���l��Q��:뇯O�k����L�zxu��d���f4�+^F��.�t/�^vX��$hbЇ��:�������Rb�=����Evܹ�#p�zT�d����|�aƩ�岞s�4��N"�HM��}?��П�wS�^����2��'�f�o"�Ok]۩$w;��r�n\��PNbfog�:ߢ6Fk��k�">�~ �*�!�q��ƨ��*���A����M�:��J��7
5҂��+�c��П��H��ЕT+�,���1y<��Df�5�a8v|���i�Y�F�v�j�����df{G�{Γ<�ᜊ���X�K��ޝ-j���Ry*߄�F$E�{h�^)��M�g��t�_�A��T$u�,cZ�J��y�t�q�=v�v�5'%�O=͞�7
�c{�ӫ����Ek:��e�����W�T�8��xiK���z.���!Q���[Gc���0�R,�������_"���*�?����
��z�k���׆)8O4��m��&��ڏlUj>>�/��7.�lTf"�eEC!m:Q�;H�|u�1s��+��o�^Y:�8�:���A�v�	�f_�g��V c�j�Q3`�XĻZ�6n�3Ch`T2�O��Um�1��b�"f�Ӆ��K�S�k���N=�z�e��ɽ��Zp�6
0Io����V��s�����E������+��b3dt"o�$���ܲ2,>< ��{p���:��lW��� �"�htoaY7���F��Okg�4����?G�?����L����� �