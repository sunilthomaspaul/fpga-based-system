XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���A��Ζ�S�éMDX��B�,3��ʽ�N(�����Hc���|�Ŷ�6O�{���x��Q���s��sǙ��~���OXtz�+����f#���'������U�vk�A�z��@�o�d�����^��?�K�_2���,]3�U��8繖8�
�9��-��GY��4������lq����#\]oB�p|�MQDS��P��e�WӒ��̧���NF�a���>�vB	W쥳����L3��6��kU҆����uUo<�ih�Ca��Q��5��a��*O��Z���-[α��[�jfc�~�e&��%vCJ��ֆ$0�[wPI��@$LM5ʹO�n�)!�����Ax��8]cGΈ��T���v�o�P��_s�D��^��$�㪥��U�z�����Y/��~h`Ō�g\9^�����Z
�W�l����7i�30BF��;�gb�G��I�����X��kx���	���!�|�w�3c�I�y��pk��v�E���Q �>Dx�F�L�-G�uV׏��v�����
�N͵������H@���*
��{�`��gg��~�c}���3O�tNa�d�a�\5��N�����t�3O�p�G��i.���׹������[�xǾ����RE��� �,7��2x�c��Vip��Eؓ�d��>bSA����	��u���G	�T�c���}�ײㆥR&��գ7��5�9GP�3�M��f+�a-�,B��2�s51<��ً_�x��Hj\�� nXlxVHYEB    bd1a    1920�!|R��P�G���߽��
�y�����4 j���_O=�ş��M ���KD��L�=��V�E�Үж򹏈���ՖF��LJV��axK�M>��6�3_�E�� ������oG�s�I�=^�/({h5���d|��9��P'Ւ�K�uh���mS�}^�����d�hN~����;[9���$�:�6�[Qog�>�5�%��9�Qç+�ħ�Z��c�f}�q��H
��O(>����%c��e[�߲>����,2�Ȫ̓GjHĔ��ߒ�f�߿���9��2!�=lIe���Fz񶉯Z�7�8��H�H����"
 �u������"c`O����@�;��L���N�V�F�J��������9s�О����P�N#�GUQn�m�<V���޾��}��s&�A����.Q'a����xR�����t�h�
F��t�� �{kf�B�vny�N��*<Y�ٟ�>i�l>�x�u+�Ȁ��#��7��K� �`������_��'����"��?x�$+���4ؔϨ\������X_̱�&~��r��6��J�P��hx=A�I�W�rN����	}�5�pP�4Y}�<��O�c	9�t
��h:�3K�}����M����Z�X@�����K���yV�v��3�'�[�'��E�d�aA9Z`��(n"�H���A=��m1��=K1-t��#�E��"�����2aY�	�����U��m���G�:�����������8�4*�k�]M�X5:w_0���fb$	��WxE�k��\�'��3lu�-7������˫?@Q�Mr�=V����x���Y��$����2'=�F;.�?pY�̕�Ԁ���	[޻UL'�ܒ����u^ؠ���y�Q_�E�-��튓"�-q�LOq.��%Q���$�g���>����.5u6������8�m��Mvh���=>1)K�$D;��n}�$�<++ϩU 
��)6�؏����)ѳ%o<}{^O��~C|gT�)��j>�R%��F%R��ԟ)��0�o8���k����(��� �����7���)��SN���x3΂�p��_9�h�����m�q��76
\J��k��d�#�M����<5��A9�ӂ˃������JP1{Y"���aq5�kK"�0�jw�Ep��{��n���-���#*�����32�v�*=;�r���m�%v�n>�	1���I�{if�.��#}&k`�x�J��Q�-���uO
�P~��R��x&����̓����$g,��.�Tn��Z��x(6���$KF,D�'� �m�ن|���` 3��V��B�Q���JT���b�$��'�A�C�f�"WO��Vd�7�p[MYm��,�h����*��5���d���D��Jsb��H㷥����%�����/�����	;�S��8�U�^%���X�R�O--�F>?�2I\���R��1QV�(��Q0�]��&[�`�>Ԯ{�����:A,��8�eT^	�a-D���Y/}6��a�2�3!�+��ud�P��Au�k��V]��L���܍"C�������c?u��<��!7@�x�Ÿ<+lʚ���8�5 �Bؑ�?��ܨqv�l��'@j&����S'��y���_�X$�6��۠1��Q}��oշ.�xyn�+�d���ߘP TN�l�I<���!k����}R�J)���,���L�
pų�a_� ��j�� m����\�w,�Zp5G$�40���H@�.]�c����{h`�Е�e����|?7{:�3p{{��%иZYui}.���-lG��ϑr�Or aU�(%d��/�&+q2�|�/�"dM���h�2z�`ت�a5%{�҉���Ƶ�?��L�X��3�f1j3����v\�������t�T�+xъ�>5rgb�}u�'zE*�,�Ű����.�ʊW�x��w����l{4P�ٓv��F7g�:�t�ۖJ�6��\q��T�/�ݕO1�c�cg�t���t�޿��cʐD��q��iI�I�X1V�#�ԣ��������P�t�������젮�;u�u[$5�w:� '��g%��g��la��fF���!)�+������{��!p��)ճl����w�����������B3ޱ�uΎۀh�e�n3�ng�Y�@aE�y�n$��`�S��v�:.1�SS3��7�4БG��Ra��;��Gi��pP��H�m��'�`�C�%�Y�}M������3�7ukph߻�s}��n���5��r�r`���;D;+H��		� O�!e�K�.��?��:6K��3�w;��P��{e0���~5&=�rҹ9 X�_���1�9�WD�h�vN}N,(�f�~�zV�\���/�)}�X����t�uS0cT�$ʛO�Ѯ��1|dSM(^���%'��B���߈S�-H}X��5c��]nɬ�=zr(\�׸.w�Vه��N��$�Z��@�eɁ��W�f�.��/�N:Ѓ%�l{��\Ph�o��Т"\���Ga���en��NM�O��>N)�}_/<�4©I��W�q�%����'F�t}���Y���+ Z��ɏr�H����PK5�ݧ%�t�@кU�5W�=J�B9e5���(�N	'ډ��F���z�1�b�C�N��
��υ�_2��9=�i�C�G΀��k�y�Z����W��l�Ѻ�U��S�/��ݬ8F.�-2���b���ٵ��\�Ln�I�/6�ݸ�{���O5��þۨZ�X�Q9���2�}	�/8�|)9���koe�y��	K����p�/ϥ�֜�7<qs$eN���M&�a	Ɛ�k�/�Ct�,�r�� &+�؏2�2ٝ�o<~NznO�n�w��s� ���3ً�(��}��l���3������x7������e��F�~�;,� F�Х�0n]�G12�����;����xy_.�%�tO�Ĥn(U�����K��5f�
?�yH�����lz�M�ϔS7���E]�>+�����zJ�`���'�G3|���j.\�o-�D ��okd8ߘ�vt��!���S��iH��Qv=A
�'j��>p8X����}�O�����@Щ�̴S�.�6��72��^#��G�����4�C��;qp������D����(E*#��%;�r29�_��U,n�l�I�����{R�	��t'��A@!6O�8�d�(��U�񼎈��(*�Y�<�k��Yb�+%����:�� �����E���ͥ+�®�E
�Ε�wTa~	_y��m��o��O#|t^�9�l���]~(��א�'T)3&<�%hpl�n��9�\��Y�%TX�N�:C�,`wK8�*�7c"��ʊ��Õ��e��u���@/������ �<@*�1�X���|�mw�i��Ԧ��91�QĀ�M�F�eߢ�D�%���C�z���D2Y{O��^�2p�l�#z�'Wd�4 r��r�`� ��v�G=�F@����� U Q4�pK��~���>X��e|d����}@����[���q�|%M�~w�L��3[�bv�d�Ju�$�ʟ�[d[_�*�ܰ����u_`����C�r�[&��s���&�Sjl��� @��>8�{�ԐMT��"�c�Xw�����"��h
yM�A+�bmb�_�}�eb�̛;�zQ:!&��ccm��!`��St�����9 ݶ�;��۳�OY�%�taZ�b���Ko��|�ߩ��m˺FQ-��^�U�5�"O%ҧ�ћx�>Л�$�,L����[�LZ���
���3�ݮ�q��{{1ܖQ�T�{��m*�=��`��=b�֥UeY�p��Hh�pe�K��޼�5���b�"���1��1���/8l��}�m�Y^kW�����Vy|��Gl�T�`�3�ͧ��QϾ�T�3_p �f9��E�	�}(�]�M�\R����!H��9P884&�ǯ��KI���{���	CH�������ܬ��;��s������i^HM΀� V�}�6�wG��OJ�V�~�pO,�"P;
�D�W)�. {���[l=p��l�jlP�Za,ˁ®�J`N�A�:���n��<�y^_��_��c���+dq�٤Y?ЀjP���ΡC����P��;<�������|~#֠&*?c�v��ȇ�{���[�R��3d_7��`W�Y1������
��rOΐ$_+~��"Dg,$w�mBt�"S�����~|["Gp�,���3��g	��Tc}�@k�-��RKa���G���)�'N�$Amsz;�����Aѣ�$}Q��b���'����ٌ�VV�3��N�'���[����^)�{��
P�0�磯�I,��������F�u�d(�I}9>$�X�[�{��@/mb�qG��FH���n�.!���B�%i����cqk��@wG��	���)hrK��@NN���S�������؋�=G�n؄�\����-]	�O��?Ƣ%��/���(�U6��*�mֽ�Fy����)�%�IE�Q������[�8Z;k(|��D������N�5���}+8jf}e�FP�}�����^R�\lI�C6|������j����!�L2�i��d�c<�sP�i�w���h
͢��=�r	����[��h�n�Z�{�i�a��Ω'+�k�JSqJ~��,����-^I�e��]��w��@�l�+��3{!��Pm �۹8��	!	H�m6%"��Ws�A�͝�����u����JXgp�-��
�T�m�)�Bb��A��O�5����;��1�N�о��C動yod.�ˤ:�OU�z��V��CȞ�&D1��\��R���h.���WN!Cl�o�,`K�{K<;L#M�/,��m��z/Lrt�4˨fA���p魦���76}�nf�h�Գ���e�p�ۃ�̸B�5��3��@Ԇ���<�dH�r.痴���=�.����U%B�DLp��yD��}�?�!�(�E�$T�O��a�$��\P�BBѽ	i'�ƃ�9'���tL��G�] �Tt��?S&�����[17S�q(ȐL�c>�,Ω# ǟ;)�U12;�a>X�j�+�(�"l������iȼ��]Mbu}��d�� t��O��䌙����*�H�3�a���k�@�Y�����P��i�� ���x���۫���Y�'�)��$���¾K��d�ӑ"n���+�?���M��+��k�a��	��R4�xBb��tҍE�����fG�+�m�ѐ������R��ӂ��F�k�:�k�m�}4o�U��	�o�����:{$ ��{�
���r�fK}Jh3�;%�mN���*��a3�C3|Ҝ\NL���jk�f�#�@���5�rbo�l�*\`8h�&��1e�DL��zQ�=�1[�@�
' �j�7VIn�GAfq
�Ƈe'�Se�+I��Xӓ�Ғ��m<����ˀ��2q)�UC��sN��S��T8���[�)<�
Bb�2��J��]�02l�������DF��� jc�5���C{�� ���G��7H��WGg�M���Y@��$M��ޜ��.���
�lVUGxd«���-�!�jpb<�K� �z�}[e~��ބ�K�W�If��핿�>,�sY�яA�txb��u���w�;
�M4
  ��<}�&C��:�E�K|俒�Z���80S�ۑGw�2@���2��1�*;�T��e�O)ﰖ*?��h½4�A(�_�$	-�����Pj�"ڱp[G�u���2Y��[���i?���|�#83|x
�ߺ��k��0��|���N�~#7󁇓��[��%�I�ht���fP�o+�a<�L��3�����{Z����f�:��16�Fr}*�s��9�Uޠ���!�D[������_��U����!d)�`���;DH��}����)��D^R�Nl�J1R&V� ��J����X����+�?���D�'�H&�A�%eA����8���n鑖#���i�-�����9U_j�fp�a�GN�+��c��\�^�X$.NT���>pL�HB�]��xc���?�͋�}@��]mKm�
��)�pT<*A,TasO�&m���J�In�[Q�Yd�=)����%���67�&���n���V�y2 ,���HSz����7� �$}�SL�SnoRt]�4��Z(����R�ң@�:#Uui["��zIJδv�߃	��\l�:�sX�d�aɛ@P*��lZ2	Y�ho?����c{߿��.��f�f����v>;|ˋ|�x}� ��U����59Z�V��ے{�oJ�'�U,�+ 7�54o�)�����݈Bږ[�+��;