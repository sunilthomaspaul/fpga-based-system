XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��
>Gq�bQ�Ep}Q�d�r�*fFe��AJ�]�g���Q�Q�{.P����g\����� Z)y�rM�x��H�ގ�y�%Ϯ�{u�4ELWp��r8��$�|eA�������6;�5iYڲ�`J��ⁿyP��6����`/o���>0-�V�OA�fbQ��V���Q��|90�,r�K��娙ٰ�"H�Q��E�;��x0i�rTӅ} �G��!��>�&9�i����s�\~���G �|��D?d�h�D�yDLJx��!��-_���}t���k�	����MW���~��tr>�t�{�^S8rQ�Z��{9���q0[n���wE+�G=�w����&A8y��@����<4-�^72����+�I{v�����S�l1��fR��U�&��Pr'��7M>pv�d�Ǧ�+���������M�,��E�����h����<�Y�/�.���;�xE�P�nl\�kUZl���ĭ�66��� ���ڋ��h��8x��DX|�b���֧=Z���c�~Vtk���C:�KR}��Q0�%�6Al��B��*�Yo��M
g��E����G�Ac��0Ӧ�0�}?�jYgVE3��t���Ѐ���M?)X8���I�kfMH[֕��q'�t@��ge�5��kUJQ�=گvj�
�����U\��E�0��ǥ`�"�!�%�Y��xN��HXيg����Ns�2i�'���A/z92�1��n����������/��`�XlxVHYEB    38a4     d00��n��}���Sũ�e���ٍ��|��?�^�A�����@�k�QI�����'�2�4�F*}�-I%�NgZ��]umE<�������9���p�2؈m�{�I��R[ܭ�}e���>Z��n6b	��he1 ����)��:�������U��U6c���s=�!C�(���cKW��b�qY�
H�i�U�/�}�0�ӳW�I��]QUnc��OϷ��H����xFކR5+���މ-��#�g����p}��$�^��2kK�B8e��`�F+���E����Rz_��??�օ��A\d�9��u	ub��2��a�sp�>9��%F^�8��A=839â�k�t���⎿GS�S�����k�kX��o�÷������2��;�W��M��H��V��N��oe%�H��!wRk3�t<��8�(��'7�)G��g�W�?
:C4�c#J����4������Uo�ZDo �v5�3��T��:�[����0~?��	��_/l�1��T�&Z����\���{�rh;��oXt��{u��"��YM+t���^�K{!LS%����X&�O_=>n��-m��i3r�-T�7@��i*Ǒ�ǁgg��$��˺{j�CC��6Afֵ�~J.�Q��1tD�s�=@vm��3T�!W�l���&��4��RaO�tЖ,����e���]4�/r�f&��إ�֗3��L�8��w����|K��eϓ�s�|�t�t���Ŕ��Cr��G0nf�������1��6aqkJ�Q�b�Ո7�]a�L��1A#�9��]V���q��1u-�ǫ>ٖ�^0¶3`���>t�JԀ�=�]�i����F17b1����m��[�P_
T�S��`0�^�"/t�:�蕞k8�l$='�oH��g�]I����%$X����(�Y!E�g8�5��
�mP�򌚼M��Z�e �V>���*-�E�\2pKCZ$~/0��2-߬U^�>��[P˃�
�nE_Z��G�,Q}�~Of���j�;*q�a�3;z~Y�R�F�-�ǔ�v1��y�6��6bȀ��<��x�	)�#������.��[���d 0b_v�gR�x�INK��b��/�A�}�������鐴@z"����إDO��=ҁ{i���GW�I~�*���l�2_�%�l�Dx���������I<@*�7툸Ib��C2�+k�Ӆ���o(�:I�f�0�A-�Z`CZ���F�Cy9ũ��� �aXUy)�dV�<[+o��߀)5O�@���{~���GD�A��'E�Q3F��� �ltf/=i�)������<Z�x9��L wAX,�5~�⺔��lB+��s׶#"=��z�h>��Q>�&�J�Z�5M�o���'�ͽ?~e�e�z�*a�ez��>���_���ê�"p�!
��$Ȼ���C�!�&�ɻs��}ʲA�X.�fЁ��[燄�E��N�QX�Ã.Szج���	��n(Zj6l�&Xd�|k�O���0��>����/�n-�����1#��zΗڅ-}�Ȟ;`�b�jJ�a�;�E����4����u��@Lta�#w�#u�s �	�S�u�;�`4�����ғ[��$��_s��e'y�^Y����_�0���k��	z�����T|����ԙ�JY'菿�+��6���R��u;��>��|�Wxstſ�,o�	"���.�,`>����*'���-�k�Eҁ��\ ߦ�\׺�?SC�z�_�1�Sm�DɈKL���T%�&C��E����p��q(��tA��ʐ���r���U?�a.� �𗶙Ư$����תEw�w�掿��c���1eS�%C�CWP���!��o��@�@��V������ilw���tc�.QS���<D�PǪ�t�4��b����8Ɓ��b�9��V�uU
E�p���8Ɋ�aq��<�Z�6Tȫ�=��/#O|{�7QA���&I止3TÑ���h?���R����� ?�$٥U~�bK����iΫ8���M 6�}a�KА��-�څ
�ꡜ��ZQB� �*CA�t�;�808�T;`��j��ȁ!��5O��X�^�G�]��h	��4�XxX�x	4�9�B��-�ro����ݗ�0�tGĒ������(�]]����E��J=�@��8�;���mT�(o��lρ�6�~�ԍ޷�(=cՉ�@
e�7�v����E�]�W8�$����fͨ�n_;A4$�mE�<=_��.0��qZ��o����M�dP����i�_�>��P'�>V�dC�j���`G�%6%f��0����Mr���4�k4�э��Ɣ�]�%�E����5iyָ]́���1����S�홗���l�fR�/�5��\���
9�uH̵���B�>�x�ZF�*��
_bS��ۘF˳����&��Ѽ}PCV˳Fu��l�|���U
��d���
���O�9���]���`������y�3z����̒��p����-aⲴZȴ\��o(���Ύ�t;c7����'lt0���J4պ�n�h�`�����uo���ڛ]�|�{��ZF�Cm$:ކ���[���a��#3{u�ӛ�����-1�r�!e|Gc磴��5���U��0��f�P��E�;&����a�������;"�o�P����}Fo��{�8������c�p�<���sMc!A�;�%?��4�2yV���}���v$���(�|%��j�B����c��+�k
$�7z1i����X�����rȟ�e�YQ�eh��iJ����y$���H�X�h�OG�щј�Dc�J_9�f�e����KJI����E9,���U�)X��q|iV�˖�_�eEJ�]��g���1pŽ3D�����!V��:����b��x���V�B}���Cf�����k�XX�Bq8�3w=��H�4`P�� Ӟp�=:9�j��L+�ڐ(W3f�	m�o��1�T]�אY�㩻l��H��g���v�S���-�0
m��=@ ��" �m�6k�׀3����<��_9�`��b�؉=���TLBq:� �g�K}��)u�غ)���#c:u>�([u�B���7x����� ��w.�!ax�6@�F��6O����K��H�I/Um]oܷ�5���r��쀶?�t��5��ߧ��e���W���v.���C�<�;����R%n�������u���n��	 9Q�۰�Sj'��pf�c{]�[�$uѐx���ֿ����Q��σ��)ֺ�\�d