XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��A4F ͡����F�N�;	�ձTsӝTJ��
�4�x�f�|e���ʍ��A��@�.�Э ��?�LY���W.���T��[�0\a�T��
��AނΗ���<��˩)RS���Qh�=�4���z��|�V�_F��@b��S��ɇ>��ʲ��y�i\,�p"�Ȥ��C���a�:�rr�~l�}=��Zӱ@p�T�	}���)@�M���IYfM���
n-�0lE6�㮮�5�f���<�e�K��ʁq�GR��DEr�����ơ��l��,��99�?���M:��K���	
�,�B��,9_<2��]���z�YF��6�iB|���& ��x��V)��^�dχPXB0��ˀW|x��P$��Q ��΃���I�-����R����a���x���	��O��ʋ����,KAƟ��h��|ؠ�^)Gb�Im�W�W�}3򆙽��
��Z%w���
�5s00B������a�Ko49�q��R=C��p�����6�_'K�{tQ�F3uRk�2�V�d*�'~&8��c{]��hf܇EbR64Ӗ�T �wB.v�j�"���dLjB��pFpC�z/W��׭N1�Uni$�0F�?�VB��3����Q{K� =��OW�m6��N��Q���:f�~Sq���eg��"�� V_�*]ڝ����z3��y��"�x��ϳػ����Si4�����m��x��t�� c���h���/�?�m�ٯ�Hن	}w;��rXlxVHYEB    47d6    1030HF:��ڡ1�Tv�V2DV�����qE�Qˑ�"Q��0�e?�J�v
�%S��n-��<H��c��VQLi3}�&4N�v� �<\��i�׌���2����D�5�_�Mڡ�'\B N��)�#:�k΃MM��ND4�6�zݡr�hE�=��$����2��ײ�|q�j�X�bAGu�����ḅ�E0�q� Κ��3e��*ô�	��1{D����~����-\�e�0䔰�
�H��Z�/	��"`.+ɣ�#����D��. ��%E'1dy!-�$'���?z���K����?|��i�'�&qv]1����@�\,E��+��[.A��<\k�dl�"����~��i\[���Lp9茥0r�i�lsD$��[?mO��o��rLp��C{�����]uH�� �����n�5Ii���4/|vd.~�ӭ�&3�Ɩ���)Щ'-'�&���o��勋O�G��Mm6N6	fr�sn*:�A��_Z�{�lG�g������Qf���Ŭ���u\�RQ������Y"4e���y)Y��	�`��
�:f:����6a�BG��Վ�e���vk�C
Nt��^)v�4u���H5������ Mw�l��FY�#|��pG��21Qlj��z�̙g�%^V�ڀv��8n��M�`n�Do�:Roi+hG5���2�����g`���9����.j;{Q̉��M�Z�$� N�f�C�.�L�$�-a�$c�(;i^�G���cČCKh7^�`�Z����7���#�D}���=����-mn���SF���Q7�Hp}�3���x쓱��H^M���a#���8�o�i�!��k��k������:Ҍ�� ���������Ѽ�����y�p�cb�<�h���t�����Q�jZ��*�EB���_39 ��v����پ*�?,�	�m�5z�Viᷕ}^0�ݼO")�i8aj�#`Y�5�gfoԤ�5��=�{�EU
���tM��.�Pf�ּxЇW^�rb!���"d�v�	�~P!�K�<|�ٍ
P��}�w����Yi�V

j䤯@�,�G������@��Z��t;�$ܠ#�YX�<d��W�d��Am�Wq��3�|�s"x��q�т:��vˇBnZ�3��RBl:��=1h2tzL��"���Mw����A�ͤ���`7�@�G	P�t*#Eq�c1���;U��G ΁'2��%/��2U������� �N�/ ���U�>a	!L����P��~���O� v,~e��J���R�����qT)�\����T�q٠���R!g���|یm�]������1}���k�����s�1F��\j�uQ�����x}�,�V�-q�a��	P'Sɞ��hb4�a��:�u�ɝ�:�.�̽����A�_&�FJ�I��El�5Z��w�/+��/]����O�}��J�q�h2E9�:
m��vD�J�b�Kd�dA��J����1�*�9�"��9�e�/l܆&4q�b����3��Лå�?�2�.&�F����7%p ��EL4�a��
!�� ��t��/��-،n�]�p�
�Yi�2��I�m��ݽwyס �D7�ΟX�J��t/J F_��(���b�L�"A��db)����m(�#����p!��f�q ��Щ�'�?��c�[#�1��緮�%��iR�y5ggJ�~X{��$�{�ک�BXL�@�&����%c_��o���e�V�D��NnV���Dǥ`<}�?b�z�=�UHx�VEyF nKc�u:`3������0G�00$A���Dl�e3�7�Hbx5S�VD��\�����J�J%s�\ި1eN!g�c<R���T��w�#� |���|�G>���Q�ﰛ�ǧ�����`-B@�|�9��u��xgֹ*��*�#����L�#F�͓Q<��ϱ@�5 �����q�u�OUo.�hf���RQ��n��#��e?Ė�#֐3 ��d�b��˖;��r(��-�{=\���.�5����xi!P����(Ra�
�Az0�R��P��2��_��I*
��o��u�*��NR7�ejz�r���<%k�<�i"��-3�X��;J�Y{�wV2���� ���&.�Y����|�� �b����kz��}��"�
�YB`N"#�4M>��(
��ĖE���G�B�ա�f$5U���%����R,.���*7X�� �L?a�y�f����[���Ƈ�Nܵ��W(c���G�y�^;o�̒�LQQY�S�L��W �a��k넭���sTVL���6#���Ԥ�+���/y�=��6�j3�� 5�ܦ8f�a��q���^;#r7��:�F):M�5	��c�z]ʩn�-��^uF$d���v̓��_���U�P.�i�,���ʛ;z�-H�NS\�7�Es40@|F0�\m�l/�kLhvB�9��/1�3��'�]���O����;E"!Z��Nsv���g�L-�~�L�X+HJ?mS�,ʜV{kQ��$[�kc���=���;{jkz�6�����p</"g�^�}�@�^�[q����P�����~/�+Z��AG�5�l���i1�:� �*��y��V���X	
1#�<�Y\��8"O�Vm�����i%�aj��tu���=;��E��}�x�}1E�`J������S���Ԛ��"^����y�8�l8�q�a�H	nX�Z���3����L��p�Ε~�賀^\��R�W�X�N��A�K2�[8�scwKD��P
4ѭ"� ��Pd*��f=�dΣ�?ZF�ٓ�1m{��Q�YX�ObX��Bʸ��FY9�ش��Ebn_5�����}9[ �a��@�G����*���p�2*������a���U��_}o �M�Z�ħK�E%+�'��Q�?��d=]�;Į{E���?���Z���v)�
�*����D�a������E����m��M�t2�!�g%f�ld�/��q�%M��,�4��ݙ3�l��-�F9C����]@�,�'��[&x�Og�����^�2	L��ݧB����ӈס�\*᠓�1�b�E���y<x��@��8�bL�"�s^盗\e>f�	U(ݕɻ�@v��8 ��!�$}Hۺ1rhHP�)��),-��H���	�����D��ֹymrP�bi@`
���M4A)�Fs��Oj��v���jR
f�R��*z�Q����~j	i���T���w����g�PS�]Kd�[^a�
����|�_�����٣ԫ�7���Ф�Ө�eE�5��ĝ2!�a��{�_i��S��z�ǡ)��)�3x��V\w��ܗ�����B��|�7%>̝�0����1^��k���8HZ��Q2��SF�ѮLT~��9؀mP��4��+��%0����S7P,^$��x,!�����_ �eÁ<�ʷ�M�7�oK��	�ۗ����J*���Iz�
���N�Dg�#ވ�ݕ��3ny���ܢQqJ�<?�䓥�ҭ�t`]��=�J�W(M������ؿ�
�X�Y��'ָll�N��xB��a��vzν�wx���� O�G��)s]@8}>ф���ZV���Kstj�Q'WYt�I��;����cA�k��R�g�=��/5�u|�bǋz��P��n��I���MM��U�р���撁�!넜���E�ж�5g�r�M�~�Mo���o��$��/����n��2׺�s���`Y�;
��W�&PQ��l^�E��0����>����K+xe��+�290������ɬ�0���Ԗ%Ǆb��&9�s�w���$�� �	n2y���t6p�ө]�B��E1��@:�����7T���z|:	u�����6Z9¼��Q��!rv�%ϕ�;AϷU37Nhr���+l~ߏ�(�-�Y�P����H�9D�����i�߾9�ö#���NZ
�tJ"�𓪉����Lf�������8�N����t�e�"��ǚ;?��$R`�mQ�Za�er�'v�Z���)]�	ͤ5B�zObo՞0�+�� ������*�rҫ1t@V�x��G�?1���P/�[�����2��"��i�<7�����,��ٓ�5���s�