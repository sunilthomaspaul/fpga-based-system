XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����S`k\�x���QE���2��(�=��`q������s��"�[�ފ�G�lAhk�3jl'�<����X��2���:X&�r�6&=�
���=#OἼYc���&�����؉R{:E��I�I�' y��]����=̀$i<9��<|]'��`'i=�Ka�M���(;���e�e]
ݰ�GD^������5!w��#˱��%�R�|�W1v��.w�vEA��)�kJ�U�r�;<����B��O.?�L+��ʢ�0�u*�<�0�����%�A�x���^�y�p�J�m� ���9���ׁ�$�t��D�笥��0(߯��W;
�����2�"��h�:�y8r*����!~U��ֈH��C���.�m���Y�:�6�C���#HbB��N��z�6�ɮHb2������ttI�JEhg�	��$���q���&�J�.��k�
���3ZF^3�Q���c�,V���]�Tu%hT	Q�c:rmVag*�5��K�����h�%֓X��/>H�z�r�����ɛ��<u�l���=�EDqI�+v<*���W�~�̣��������:4;��> 8*�ca?(�֤/��=j	��NFfo�P���
֖)'��Q�Z��W*�<P��iAu��ԡ:�m⹨4�X�Q�ɼv6�f�x���uG3͌�m�0kLG�?O��֑0]b�ڇ��j��!lK����Jq���.bc.���F��S���U��l׷G�ԋr�A���?.�[XlxVHYEB    4548    10a0��-?&��nr���/P���'h�Lzz|�Q�����|����|��Ӷ�3�v�uB!h���*BY�BO��=�M0-��\-$��z&�{=��jN�+?[��ց@����D#=ajo O>P�� ��[q[l�J��w��_%"������t�=�5�J�(Ӱ�B
 �C!P��X#sE�uYϒ���]T����q�&{o�h.�
5�`�{DO��4��4�T��D�J�&yi��F]LIq�	�����nj��+^[��\�`�tF�1���p�Z6^�gȶ0Wڕ(���K4�f�qI�J��%)b�W��0r�of�������e�L�㰋����*�(%��A%S�	ђF!Vwz�~8(��W�/�cT����]w�c��𬄱 )y"Ӕ��٨������$���*��<�÷����|T/�_Qf��)-"��r����&N��Q�~�Pla����1�;an�|�Ɨ�H�
p��-:��w��U��v����\9Uo�<S�~�����ו�|8ѯ_��4��Q�eL��E�b1 �Κ�����4�%XN���C���9��z<i�]�RK	+��*�����j��uRC�ڸ��l.ߦ��@~�&���se���+O�6�1�1V�p�^�7�'��E�ZciM�ws�~``ᆲ
�����2I��L���J=co��'�����n��	�T�Qۛ����&�'�6��X���0�bc� ;�9	iK4;�xɌ�
���7�E�6��w�0Eu�� ���}q�R2;�)�4T��C{s����)�2l%k�Dл�N3x^�fSI^�|��9`a(
��7��e�ƀXSMsd��h+�q;�xY%�/��M�Y��b�s���@73ݴs�Q4������s��8z���PlCc�by7�_(Kc!�����̥Nܬ�M<;#iK;~��a{$^����j�n��Ow���+����s��T�3D��}����R��#�-��1��+�]>'{��.vq\rdz��G1I4���UDս����y��[��ܧ���#�Le�f���f_8�. ؖ��R�?���c\k91��3~�r!ʳ�G�!#�������{<#�(��u�1�V�=�����o��f��^כ^yn����W1?$�[hh,f�WpP!�ϓ*�9�I�L�l=�q�I�-H?�j�Ğ%```:R­�Ik$G��cƎ��M	�(�hE�?�M�Ǟ/�_n=��q9\��ɟ\�UN�ϧF��ڿ�#����
S��;���ͭ��QGb��g����/�15v��g���M�@tTΑ5��������R�	2��GW^��Uj2��<���fYy����E(��ÀDj�33$c ���R,g~��h��Z�+`���N+ׄay���ú�hH:�V
V�#�gg�D"vT�2?����Z�#�y�E��8䊖G���߸�v��=σ�:򌒵�����GG�^OuS�i�\��������v4����MY����+���zf�in�̌����.X���'�<�|ϰg Lށ^�-����4�m�~���W2��x�tzڬj4z"1�]�Z��C�C&̍�2􇐃FKҸ�k�Dm9'u�%����R�M!x���v>� Ž�/D����@f�రaCPP;k�/���>��� �5ªb�H�+4Zv'�ò��*l>�O��>�,��������+ݿ{P��W��� T)Q夦^���b�O��0�8ea�A�bS�@4n���)�m逦��ye�������aX8�k�l|7ݘ��31�j
�x�`�5f��y�a������V���2�ir�s@�݈�[a�'z�3��5iSq�Kd7?`�q����JHY��g�L�Ͼ��IN/�t��-��^혤����
���8g-zco��Ln�o�S\��[#O�:q�~o�߿�NC)�lb��l�,�E�wjD�;�#�v�+lǲ�J9N��3�~��:L/�����. �<�� �&�'I|bϝM��_Uܜ�,�NL���j����HW첼�����4�C�"�S�C�A���Db�0���|�۱�}]3s�To��ۤ ����G;�kq�<�o
�׌<N��Yq�qMR�1�-6��"����	'�57a^2"Uzl_��ֳ�1�KG~a%]��חv���jܸ(�ㅤ���.��2����æz�'p�+V�)lɉW� h��`�C>=�yG��*�gڅ�.��i�uᐮ4��FUT9��!����YXK��:N'�7s(/2��y���j�H+������.r��l� K7�Z�	��^��
�ܳ�Ԇ�@ă�D�1Z��tP�Z�:/1@����� #.��IWS{Q[�H{mL_��`ᇊ0����U����9�F����SxN�ܐ�3�������M���)�\�gz�� �3U��nM�`,�h��P���+�œ��;�k�t�
��Q�����|�:u���9��]<��X��`��
�6�*Cl��;��'"Nڹ��O�ɱ��] 	�i��f��=�V�j`[��b#����ը��y�s���MU�%΂K'�0��+�~���6yoq��6�w-+ q�]	��-��]hF��zxl5@�}֦?@���N 緼���!�,�� zμ��D͝��*�[�3ګ�[Bڥ����cjNKZ�a���k���/�0n�p�4�T��偑��[Sx�ޜϴ�4�e'�o
f)#fx��L]*,wD��j��ֆy��6~��D������]��a��Xc��BX�s�o�t.3� w-����V8�c���_
�C�����Ú'��~sBC|�S1�Cس@x�C��D�O�",����1�5�HO��ז.U�ч���艴�u����c���C��7I�<�륻�;?���l�F;<'2��j)���GQ䞕J�`B�&���3��
qx���#/����
��C�"�|:��/���w�����G;0~;��µ5���|�l(�(0��i��h�j�=��N"��n��IxN�6��H��{�7#(sLC��

4�`��uO�g���� ����&���DQ}�h�W�9�oøn�L8�feQ�?-Iع8��M����~�VIK�)&6�-j|.�$'�ކSKi%;�X��Ğ
9��N� �e��&WǌDǚlс����)���6�)|?#(�a����4�O?_��w���-S8�P<���q��-L�N�f^A���u�-�j����CV�O/ �hX�4k;��p�z�����a�k�y5:���Kʎ/V���c�p`�Q�Р �t��)+����,0��{�)�Ic�W�Y����	���@�zD�#9�Md�>�GhfO^�c�Wǂό :{tt}s��!l;o�*�)�G�yJ?bmdqi�t�@�:���e�Yӓ�N�@y�W��&��	#�Σ(��&�?��o;ߏ�1 �P�]�^�¾���\F����N`IB����>T���,̖��yC(�t�H�A��Rq`��:�ޮ;C��ԷI�2Z�������ζ$l��堘s폢���ҵ}1�c�V�-�:��>>R��u0��=V�[�����8=]"p,��eN�4�,^���g�aL�J���������e|+��&n��	0�������/7s��%�|��:�&R��nTm�X��lp|���	T.�?oC��S�LA�C�ɂ_ �S�{ƫ��HE��"�'�2uP�k �b;QA�����[@���Y&���5���Vl�l�Z�du��wF�L��n`bC����	Fw��>����]#mP���Mrlw�=�~�� L[�I����ʺ��j��ru{%C4Rh������vo���亓;aP�$�Z;D�t������Ul����/CzP�D�(�rV2�D�κ��� ɯ7�4o ��A����ȁ7d�d���W�[�ﱑI0��� T�����Z[�U��Q7�H)�=S~���y����糣�y���������`� A��j4�u&́\�,E;�mJ9Lm�J�\/��A�06?���{�d�������;`9�k�ҵ�)�J�Y�J�
?>,w2wv�`s�'�ƿ�Z��\��$�L�^��� s�;w-#e�Q	�%��+��g�A��v����"1���mtEw��I�`v��!����!�Į�
{x��������L;�`���C`�׬_�IB�bny�<�t