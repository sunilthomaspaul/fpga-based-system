XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����+%m%�W$]�C���Ϡ6h�_v�js���"�q������
��s&�i5P����*3�6�+�)f�����˯�j��꿱C�Y�&ʭ<� W��<뇝4&��F_ql,XJW�v?�Z9kRh��$��ueKQ駉o����u���c��ԟ�`VF@��s�Iw"��R�DECC|d��9䅃|��jX�BQZ���.OiÒ��"u> KF��X	� ��X��G��G��M2�YsGM���Dt(7�Q�ɽt����r�����I��w����2�6�,�	�B�4=��!p������&�m��?<�I��Tk�+��=�I(�Z������?r�(b'��:��ʌ��m���w��tx�
;�lJ�(��5� ��L�iZT�����pH>��f�}	?���p�r���:��&
�砯���CP�N)�#ؕ@�J��n�w�3b�?�I��#�D�%`�w�����1�R I�AC��T�)ȿ���Q�t���Ӹ��a��t@HJ�!.��4\`. �+����:<d�����Z�>�ȥEƊ$�׵b0WD[}�ǀ^���ļT��7T���U.���"Z�n���w���d>Dذ�}l�D'@J�IF�y%�S	آ�0�cB��d���M��N�I_p�(�r�$� B��bT��m'�/T>A,�|�.���̾$�|@L�4�S��!��I�giP�*K��QL��S���]fC�ި�	���Gt2f�~�S2��klJ���"*&�����O��XlxVHYEB    1661     760��J�R�g�e<�� �S ����}`���ޘ V�]��U@K��r,'I �%��G/t}\��.�8�x_bծ��Uk�5ÅSI%�*���?�݆_��C\T��@?)��|2��O�����d��J�&V�>'#�۷�y���7�2�����l%�N:��>=`����� �'����LG,�JH���/';:�s"1��\3Dή�ǽ���@W��r�� �F�,�Z�қ%�@Y2�GQ�����:�f�5�⨕�2���>�%����#�ǟ^% �$GԒ�D=�`~_/�+� ��9+�#����yC��=ِ9F�u� ;��U2�>�j!��:���fRZ�@��*�Z%��hbIԩ��E{�W���&>���A���>��{C���M��h���EY^O:�h8cLHkT}��p���8�T����_4�y���������Ivz�s~�o��9T��#nHÊ�ax��ֳ_c!KRr�]�c��H2c(�+�~PѨ<ƺ�<�&$6iW�ӽ~���/�p0���,EB8������p^���A�F�DP�����Y����z`ů��C&�4�������#7���1W���L��a��_�Yo��=���X����$�lLH3=OO
Un�oV~-�~�\vN�e��)�W�`s�z�	��g
[
Z[m��Ŋ���%�Ғ����uץ����^P�TD�L;���7�m�M���'(X�9��ZK���-�"![�ǰI�k�)!�i��?W��n�fv����������a}M?q*ɞXF�7;΄_bT2Cn(��S�c�ͩq?|�kn���$tz��W85�E�@�c�jWB�UHy�]x�jJ�ӎ}t��("�L�LP������0���*Uj��7��ˌv����9��S�o�~��.B�GW�`w�s!F��b0z{���OZ3\��G���Eun`���k�^1�����}��� 2�<͗�b4Ow��VoY���H�t98��+[c+�F��F��g��֑� 
�c�҂�p\���_���8�u#���t�y��rV[��Km�Rr�:���X~.� ��H������:e�U��y)n�t�H���C����x2�7n��<�׺@qǭ)42E4��� ���%H*6��#�#��$��'��l\��/V� x{6{�;2T��h/�[�A�ov���T�����@���x����Io~�A�ݕP�V����Daપ��Z�sIa�H�r��������o"�3S�bt��UOy�E����0Y�L9艂�F�)��B�-@n��{L�7�ۑK�Cz%]>v��|����|��lи���l��n�o�UP!���HKt�(;��TO�q�Ĳk��Ƕ��3�X�&�����Ԇg�@��:�1����-����?z�q=�3iSg��
�[NWR��՜t~
lؽZ	�#u?�,ڮ��ʃ�L�˴m�ws6���7c��a���$�Uh'�iFQ���s��n�������YM{t��z�#�����l{����o��Z�yk`������Y�Z�C �G�לƁ��� !P�1�;��iD��P�a�o��t�]������IsY������n[����N$u��|ɸ���ȯ�<
%�?�5�x�l}\_�����sb#�H���Ii�|l/�����s֝UM�]��r���:�m�x�q�_f٧��	��^S��-.��A�YƇ�a�������~��?֧P�=�G�]OԠE�[U��`:3�r8�	5�Xh��6�� {�kN(\l��~:�x�X��8z�En�4&��Ko�����=ӟQ:O3ܳ<m�.�{xI<m���!&�K��l3����kF�6�>=��A