XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��U8�ԗ�«&E���r��cw�k�G�K�`T1���^��[���	�D	\�H��r-�ZTV@��RQC+�F�&x6N�'4����B-������*�A�&���"��:k<�k��]�*dA�����(���UZ��9���u��CTp�`�8	^�]Jx0#�.ԧ�zq+}������I?w�W��)"����f	ܣX����#�,s�:
C�T�|��C*xI��C9��`��C��Q"���x���\��R�|'��2bo�b�9�T:�t<E�����8���
[Q�@�1���p��e��G,"H���s�/קO����j��x����6@�Qa_%)�~��U�:N���Ϲ�����}&�4 vYn6]�X��b	�������>�������;��-��MR4�x�TB���!��i}��n�|~�����~�`������\Qra\�7����`�8L���/b�{c�j�B􊆐����j(8'�7�aw��u<�D�Y��)DNi���tZxX(`ށ;=*��~�co����#��й��p:��4{jĬ�p��&%ٖ�] ��P��g�L۾�m}���$>��[Ӻ����|�a�H	@u/��bB` �(����'�u^s�q��f'���=G3�?&�7�e�mS��܁�3v��2��oӿ=o�ah1�]��v�����FuUMH��6�~ _�=�š�AOr�:�T(=���I��h3a��&8]wc�%�Ȫn��D0�<�X��Iv�Abd@������XlxVHYEB    1017     680eߵ��B�P�j��0Z:b]{�;	�B�E�nS)$�S�N��� -!�l}�h��& ���#?z�T!ǵfL4��@�/ d����-2���/=��	!^���,�&��.y���ӫti{3���F���"�i�k[K_�V�G��T��	X��y��M�� zC�ќh䌯�z؃˴��&8iM�,+rn��M��a&���̦Sb,UQ�8�?��7�`�%RgL���P�R	zm,Z�Z���CF�6B9KpHĊVKg=�!���1wlc�{+��
��@�r����9KU�79�/
I�<�V�����4�SD��9B:H�%�>��xA���-2>U�%��Vq� ޏ��`^�;	��C�����YiQ�wnB!�hH�A��E	��/-Ύ��\���9��l�%���i��`sE�-<�p#/��Í����:4G���>8��� J\u�����3���C�ր�9��}��%���ix���DE�(K6��	�NE�a!\�6� 8�1�H��'��ڶ4dp�e������j����]T�$���&���a_�5~���E;O^Rrr�������`�r&)`$���7�Ə�/�a�2K,��M�u�y�ǷK�
�~l/���k�Oc�\�hk~�
�2�����vN�f��w}pd 2Q"/i�p�I�R��T�����B�Cq��obr �]w�e+����ks���@߀��u0��{��.0��%�bZV[�a�U�6�����'sL.>W�Հ�[y_U�pk>}�E\�9-�i�r�e>]�@�v�e�P6�M���!@!| #l�2����1�r��otX�N>���I`k���N��Jm��L�?S�H�م�����cn��^�n����&O�	4��l�ĸ�#O,;����\;q0t{)��E&���[�5�3��@pv���1#j��b��Y�2�B�y���B�R�z�R����o#��e@��Yu��'�z��ER�v�Fmbd��$z����nba��@�Cl%�!;����	'��[�0�#W���9/��9�^Q�B�7�d���dcJ5~�4zvz^��\�����F\o��3s�%t/06�|֜�A���7�Z��6�;_!Q͘c�}C�k��%v�����9�(��鞲�����V��I�h�~���K3��ݐN!���B���m�����Įq��/�X�y�r)��j��n���|��� �p'������"�)#���1Ȕ�D�X%�"1���ol$��*P>*@��=Z��b'��2�ې���%1^Zu	�d ]��k�y{�~VO����%����"��^կ���U�j'���F�ncx8�b(��A���b�61���d��:_�,rT�ij�Ho'%`�t��˯���ƐI�[���;7�^����TR4�s<���Kn�R�Nq���|_�*�rȽvE����D����X~�~�Z��|�]U� �oJY������F-	y��0���U�����^�Ԣ*�Ż�Rܘ ڣ{�+
p�ѣ�ju�+{�/V�/	�[��O��C5����kp�;�Q���`l]hگ�ج�l��=)�ˎi�{���ʗ�b?�8n�?U���u/�D&���9�i��4$0ٔF��-2W������Y