XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����2L#��I	ÀMJb��;G�B4 �K��W�3�##yʍp�ԓbD���KĆ��9���O�Yu�x%|����������D�*1�����p��歝wU��N���Ѵ8Γ�6#��J�i!���3�:�V[�Wl��^��T�e���/D�:dM����n��(G�����vxi�����r�s0��tߗ�m�,+��q�
��H	>9��`��<q����O�oO?Й�������^���S"��7
��l �,8{�X]+
�.���^�h 2�@��C!�X���=P5V׶��g~�fO=h�csɤ-�¹�[�T��e�r4�T�>	=6�e�BV���Y)��l=.S��t
�(y�tˀ�+������f�~0IT��Ȭ~3�1FNm!zh�Pi����5B��3�4�ז�܃�4�2�U&�O3�1p+�α,\G�C�����JR�}��`�*�3�H��_��_�96ς�.��z�{�h�HP�9��$L�4-f"�b6���s�f���s��6���*�j�� ��W
�)������.��:�#�ar��H�y��86�L��!]�-2Y�W!`ʨ&��G5� ��8Ƥ��@��}F��Y�h2,���&�~�d�[p9���C�g��cU�ɯ���˃���E��Z]c��&��2�K~Wz43h���c�a�焙�O{�A���4&>�DbU*�pUxt��� �#��K-���$��+���^� �%�`��XlxVHYEB    2327     a90`K� �Y0e�[� �f�
^fx�� b�d�)Q<�N��!�5��P*"{:�ݪޫ�4� ����(�d��@��,�k���U3Pqڗ�V ҂��3�:�V����X�!l8��K��P׻��ІX�Y���~W'��UA�a2����,��?�����Q�$]�(P��ō�,3�X��6�|�3	r c�H?Ka�C�����jA&�q8SD���˥�(������,�� ����sN�Q�K�C�έ�r<�U^��r�ʮ��u�6j��`����������*�x��=��w�`����Fyo߮.\=M�,�7_&��U�L��M)�!I�W�\wr�w�C9�0������#bg��^�[f%6M�^��ˤj
�z��p�R�Y���*W��8�Pz�۷	Hv���,%M����?�>���or��B5Qw��}�X�x�h�٠\����ˀT_�8�3YkV� ��k؍��]��^/+�
8.B�O����dO�/�#Xs�3;V�ǛN����_:GJ�F������:����J�x����Ө���́\�p�������5
�r�MV)�EY��P܄�Vŵ2�s�P��r�����_�����1\lf��'?>*����9��'�)�2Dϫ�x�;%I��P��Q��^Bj�%{�L$c糴��D뮪�/�H���� ���^9��K�2ґ�w]����P�&��3�a#��3?�j"�g�k�|w�|Of3굺?:p��pAݒ1���SH����͌#+�Sˀ�������#�	��n��lR��Zd�:�Ŵ�� �����|�[��*6㿖���Ly��/����5�9�T�@T/��;p(�W�12b�s#�|kCE�z��K�\Q1�-�p|�<o�zX�La+y�زao�e�K�i>a9g8�=VYX[)E�w��;��4f�����O����ŋ@A����9�b>�_��r*�^(q�-i�I���Ӻ��x����eOG
J^��'����o�b�c]�YMF��!���E�߱�*5TW2�s�\F�f��E���@��%X����WJ�ڗ�VO7i��ˣ�����*��c��@~��_�tO�0أO�HW8�jZxR�+l�+z;c��T"N(��aj5�^��O`I/PC�4��9�`,Z�^��W��������=n98&����Sxր��������
�/��r��j%�n9/W(��2�>܈���F��a%M��G:W6`�U���͝��¯�J��M��?ۚJ¦␥���AiB[{^\�(��2�um&`ۏ����\�v\�׷r�]x�lFq�����$#��Q�F�m���#&�G�̃z�)l��Ϻ�J0�h��]�R�d�F�u�����T��$�A�fU>�E[��砗�@k�t#�{y))T ����J,�=>��q/$�QB�i�>�S�zҕk�9��N�Y�|�N�ݧՕX�CfIg҉{O��&²>�:��R��ě�M�k�dܣv���+��������ymuV�:�Q�����T.3M8)^����{�ܚ�������i����ˍNQs�}J����|W
��C�N����1��g�!)�
�� 2h��b�4Ƕg�	?Y�o����G1R�q02U�6�`�I��7�v��+ha�y7m�J��6�,S?�$�+E��'��_�e�2�&��]�vLR眒�޴ O���@���0��ΗQ���tiXǬ���"�нxD|���kt��U;Y�qh��/����C}�bj&��X���N�uJ���5XSG�k��,�n>���B��{��oM �:�M���[�f{�Wn�R��o  ��/@�:jIPN�=��ɿT���'���2)���V���ڙR7��ߚ�m�O^r��_����l���90��U��(�
���E,۩C�f���Ի�/�*K�dQ�㷋h�Q�G���_���h� ���M��C�K��n�%_Jw�,ie�bC�ue$K��gͥJ���0&jЕr�[7��5൏Z%A׍
g��A�T}�Bb���g����+����- ����J39��{�Ġ؆�#�7N����>���b46Ys,'��~�Pۉ�Y:�*y���2E8fjL�o��3��@�^�c�+��K�fu���0����-PP��>����m����1�e7�� �IV*@�4T'��X���l8����-�պj�87����e�RMK"&v�ur��}�ddM�ˢ�h3��OoK��(�w�g�"�-FV�] Y�``Z@��[��,�ń�����U����u��φ��m���酛�3X��EI�^�с8�`�E����*㨃-�+8k��Z�g��GCd����X��GD����Y''K�������ɝ��!$�3� ��wu�:/y���*�D�jVb��f����ot!�̐�	y�l�� 3�t�no	Gy��C��i�Qk�j�u1��G�F�
��;Aj�?����G�#"���R[I
��2ukE��*�6���������H�1A����Z�TJg��S�Pxǵ���B�Z.q�	k�1�fn�z�/8S�Q�q.]j��T���j�G�|8h��@I�����.�W0�G
�@�0憐���i0�J�'��c{��
