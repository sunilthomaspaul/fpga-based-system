XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����e�<#��	W���hNw�,���.��� *���)�al �9-t?Y!O�7�;pЬ�� R�@I
D���q��2�{���֟{��0A���`���'�O�����HL�{6ͬn~�0\�YB�(�x�jq)�Ւ�.0�nB���f�Â��('��^EG�v��M(���"/����I��ܷ^Ҧ����fD����j��\q�BE:"����2$�A���A�h���$��	
WN��g0���7�?7�`��TVД؝�gj��f!�Eq`s�C5�9��د0D<	H5��H�}���D�S���V��kx���N�Xg�l��4�Gv�]z��4=%��	�P^e԰%=������[��m�c��"�M������@�\5#���^�Ѷ"�����*�> ����g����5�r�LK]Ս|�50��a�����LI*c�}JiB7����]�>�����Y���eRh�\p�
�ME<ڷ����͡�$tp.��w�����k�Qy#G�8����$���������3f�0�X�T�PX��� �)�82�"?�%�Q��b�OȰ��Rڙ�l-�d�K}�N���_X}�9�9��}g�F�,���΂��D���Xc��p�U��0��!b(q�������� MH��	�L(��x�[K\�IJHn�ۗ�f2�I'�y��T�B��K�����mX�ԛ��X��7��Mp"sa�d�&;�h����hUA۰[fW��9M@��rKR�Ck�f�AJ@�#�XlxVHYEB    3292     b80���f�\xڊJv0)�D_8P����P%g��^�R����oߧ\ȞH(էĩ�g6�}��f�~f�We ֘�1,��?���nSN�I�R��0����ý)}��i�3���|]�pV�3�XY��$�t�E�A�E1M��+�yʾ�Ǐ7�m��)U�E�P����N?p�{�˾�y��;@0.� `c\��D��v���#`�p�U#����t|��UG��}�Y�n�&����` /,��n�BH��&(¿���ϽNv�ρp������
�3N�ǝ���}�7ol*�H�.DcA�V��9�3W8݉����'m��q�Q\~#���B=��y�/ˉT��6��Qm�/�xyޜv�IO���y�mbޗ�۸�c��}Cj��k�V��8�A�Z#�"��m����>��I�����Hc��=�!1>�3�h�̲ET��1G�s�e�����n$Ի��=���� P�����S�z0&
�fc�=�w~�Z��@q�/�S�jw<�\�@�L� o�&�2�_�=7�C�@��<�����`�څ�@�.�f؍۪#�5fj���R���tj��i�a�[���"hz�����V����{��%���@��	_�R�������ǵ��!"���1�����b�XӞ��iQq�t�4H��,e�D:�s�����sX�o�D5&rGc������	{�R�3=����zk���n�t������Z+"����!�R�@���K�*��!������"Xr�a%Iᙧ�$�̯�|[l���U3/�����/��Uf���������j�d�",_X��y�D�_^���P	3�<X_��U��%�����hY.��`�	������Q��݋��+���RH� �~�_�/�l9u�?�����5�Q�Tׂ��S
�ؾp
��:0)l��k�BT��o�~
��9|��<�͙w
x�'�����K�����H)��!-�� G�;br�Q�2&�-޾��=�S�Q��5��<�iІ�1��_)����>�%c���{�/��qTχ������C�;t|\eXm(����h��~�)��S��L�z���`��EK�`q|�lLGߝe�{���T���D�I׊W<)HRt���+K�6.�~l��k�q���~]���67�ﶜ��
���Q���6�$$�����{�r+��t��d�.Ծ��k70H�
$����_�,CG��aw2�ZN��ٯ�� �p7�q�o���I�e��I�#b�3�Ϲ6�� B����Ù5��hw>l6$�6d+!S�CU�Sf��[g���_/���[�+��%��;�@�Maґ>�$����FPG,	"NR�r�I�ٿ~��?�����4�7�ћ.�2�[$]�@[f��z��'�ϭ�/�L�I�GO��D�a�4|V>�%@��w���J��[g,���}sz'&��-DaY̳�NS�>�l���|{�l����,ɧ1���[k�3�]��T/�xb�����\��Yԓ��쮖R����r!g�,i�����p���z��2 ��(z�t�����/A!�J<�RZ-薏��aE^i���n�(F��)��Ka�9s�2>������d�O�hk-��m��\�Fe��� "q�ߏ0�W�1R5��B�q�c��L�^3M����Z@O-f`7��]�S�-��Î�K�^�I`��dI:�/U[���Y�b���,�+kb� ��
��$W�iL�8jȥ��R��O�A�!D���	� Ҽ |=�H�wHi¿�֫b�fF���@&��I-�qǙ^�W��އG�r���D�cR%8>�K��f��0ǆ�֛���>z���3qN����ob
e�e�� �_�oJ�CH}�4��ש�y	�S�iط|�N?)���*��8P*m/3�I*�~��U7V�#��f�.>�(���~����|K��R
����[�}*&t%}�(G�i�[̆6�]�Uǜr'�_�������M�x��I�T4z(�G�o�#��@uD���I�>�`��lr��ȳY�����s�"ܑ:�j��x���9�&�_&��g�-�y��ku9��X��(��8T-��N /�A^-���@^����늃�W��E���r�V�B0�):��,$R?c�)��F9���^�K�_�������3z�L��4#�w��:{x���[?U+]��x���D�08��񙹷aIJ/�i�{
�+���@`s/�L&�����H�!�I�|��]�@Np�k�QI��19��0H�=\,0�����à���F�.�Sb��f���i���s�3�#Э�|'��(�f��� � 8}eU7�3�|A��=�A=�M�SV%WBpH<E�� c�h	���@Ͳ�%�XG��R=�qw���M�Y�)��s0����`������?l6�ĥX�n�x�>`���8�6�sW�/Ӆ���C�D�������7�j�kF��������?)�7J�fiσαK(��=OL��Q��aw�D��\���U�A���,�9͓ #����B�#(�ƃ��o�W�E�oob�ߢ��F�-�Ĝ�N��<h�}�O<�q~^[h[)7iۥ�����F�n.����6�>1���#֮��3�[�k�W�}��X��7���v�op�����C&��?�R����N�XrAV����"@n��w{�Jm��U-:��s�dġ=J��}TP�l肉���h,��5����^�k{��kjۙ $.X���t�{��K۽��t���Mj&��<]�H<��(@z��_�e���<��si�c@	�|�44u�2'�O�=(����A��s��n��gT	�xٙ�y��� ����m�1PÏ��YK��f�*!䰆F�mTx���{