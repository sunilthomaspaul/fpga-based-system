XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�������3���Y��?�x
�����{3�鶚� S�kf��S�~꼑�U)'㻀]�`�
�����{;$��@wM� =�u?ɮc���)��E��:�qЭ,�8ύ��f_�E:!ʩ�1�{���J�Z"��^s}b�ɕ�,��}:�O�4.uL ��gy��|��G�	-G�#�!|�:�2P�C��la���&I紪' HGÆ>�AJ�:�γ��=���0���<��0�r�����EpRE��2���%rJC�J�������%����m����%�U�xXqB��6�YObt$J�Z`����cf������À�g����Ľ�8��0��<ͼ���t��������KC���iO���<uxi�a�g��`j4K�7��Tk����%�{�������s���s.�>X���~�A�mg&U^���9u���|�2H�yb2�� ]�-{F��#<�����0y
<b��9����:�8�xP�IТ���$��w`a�����]��\��%�d�gw���r�'s������6Z�T����-.�T4��Z��|]ڐ7qYӿ̼�F����X:t���f�x#�c�UPϬ���7��������0�k���d�p?n�%S��;�D{@
�k�(�5�[����c��R�DndǥO2P��Ͻ� �4m����r�}��ʹf"����m��}X����E�������Q= ���KC.G�?�e1�U��ENq��!�螬��^I�_���bH�XlxVHYEB    3f19     db0���Ϯ������h9op��q���J���wB�3�߉=
u6?��dUb?�e�aۛ%V��.��y�,�X/~i*�ӌ9T�Hd�JX��@$�{p��p�aF����<�C���i}�0C�̑����Q|R�%�D�
9A}S��(�c���Hu��p���q�K��Y�grQ�'}�]��l�<+�����
o�m��쇵[�n�r���Z�ԧ��$�mDz?�R�!�x^�N*��-�7�x_�=��]/�d��H('��}�q,H��H`����I�q}F�s~�3s˥k��
D�",�VS��6l3l	�*4��N՘�扤A����+?sW�������Z"'�)�9#�핚�moS����
�$Z�L�����Ţ(e����jlćD�5���!+�ex�N$v4��8�+����[&��&�;7���������=Bպ���P�إ����}hx׫�JS�%���"^f�s���i/� ���U�67`"�\%�ڔ�{��1�R
�[V���0x(��� RN0&R���n`����z���^����&��h�^z�x�u�֣*A�z�^�1�?��شQ�	b�	��F��6��(92ȻU�FԘFܦtK>��eZ���K �@�螔{nB��U��;��S���k�u0�l�_�����Po���|ZV��fg��*��z=�/���`�>�����)����L��p1�*���mxa�5.>�ј&a抅]��ѕ���@ܨKCw*��^�Y�6L>�R]�dW m �kv.eg->3�rl�����4�}��z�z�@�����y��M�|�h�i�ʆ�F|����C�_�y�U(����r�FF�����v�Kb�5���J��G#���HKI	8�k*,�X.���i��(�f<��d����j�N}<pR�y��v�[�}�:
8��U����mlT��.\���yg�gms�p$�i���ğ��I\���B�п����)�FİHw0��q������<RAD��i|���\q�'���b�pV��&���;bMt�d��u<r��������<"l�i ���� 6~|�h�� h�\�4�_�����vX��(i^Gunq��FSX5��� �(P7�H�+�:` 3fQ*u���*pBH(cX#�N�C��ܨ-P�C��L�	�+�5hk�1jR�`5��x��b�pMԵ=���V)<�@eu�������$T4QoҰ5�5�,G�Z7�(�|��&���q�i:_c��x�����W�l��,>ע�T�?�x�|��!��w��e6�����3�x"���;��se)d�q����ٞV �7Ki����9D�������RI�=���BR�k#�݁NR�rl�@�!dIV�B:��K����K�� -�$	���]��}n��1�o�1���j�+�J�����Q�O����%�ׂD����_��;Č�U?��q�Ox�Cj4���g�X�Es�?����qB�՟2;�\NĿ�G��%-��	�j�M.�����׽��`���{Ġ�K|V�����}�0��A'������֧��u%���݀�Be��9*�I_Kgzz]��ԌN�M�Ȧw��؄,���Cqc�zB���(���*<d|��o"wVd�n���lt�����c�M�Փ����y�Y1kV��
���*L��%���iHƪL��`�ݪk��9�����  ��;D��ľP���`��څ�s�t�u�j�YZd����7�ҔȪ9�&y�k�S}�����y���25��D��bY�X*�%C(���zdl��e*�;�!�
�r�v������<t���Xn��(ɟ�N�A��m~,_z��B����\����80�v�4>/���/�kǮ��'��o�;�~\��x���*���&qz�
`��}Ҩ�0U�7|��G�3��8%��,{����ÿ��_(���e���!}bU�t��k�=VOi�ќ�}Y0ض�v=D燢\1`�b��6��4�< ���3�"�?��TaeCP�D�܇e���j8%�:uR"��.�l�IzA�&£51�� ʃ��
�57�}��ɫ�@�(�5�b���F��/�R�/��bI����,3g�����`@��y����������R�nI/q�"����#�;���۩�I����z%���a�km	=�g�������2&�.�B���~��?3d
����2߉�������Iw�H����>-Μ�e�|��e�{�Y�,$�9�M_����t� �ݰdOG��l��f��c�ѓ�Fl�q�Y��M`{�"V���>���^����_��
�ǐ	��g?y[a2�Xh�'CJ��f,��"v�)'��L�R\i6"�Q�a���hkB b�h-2-[P�7����8�%
VR�t�7g��D!ڒZ��������8��R��� R���@���o���X˒C˕��K,���d��#e��4ʉR����)~f�{��bB����O ��<1���d % ^&�+���@	m#�	m^�cq*�$�f�/�����S��'��ڕ"���{����fH�]�7$���L��#$]O�fN`��]�������e� m��n�Z,�	�?�"׭d1䊃#��"�tט�3���A�t2��X�s1���@��"��s8��*���K�A�@�k�:���(�)���GU�">_�Mڭ��BL},�ڣ�er|����cC�GY�ҁg��?o=Cd�h ��?��y���O�q�m�p/�*�Ng<n�6[�(�F��WC�V�{0�q����u��7��ea.M�ޝ<@<JѶ^Oh56Q HB��1�r����K�+^��JRܩ�`��`�_�* L�q��J(#OyE��Uh��Ԑ����ZG8�޽٨
�wh��?3f��ʞ��P�y�{֒��(���&���KB� ��|G��Z;|���4�h�wj��� ?���������1�냦t��'�h'X���L�� QR;�48�I��YAhILy�ӯ��q��#7\Ֆ�,�����+}Rk)<?�-(n;ZoU�n���u���K��E��&��G"��˧"�0o{+u,[c�
�%Ht�&��=��[���6?7���t�§�����۷?�@k���f_A.Q�ܯ��>�5�]�.�u�9{0��'w5�<��,���
b)��TݑL&"B�1z�i\]��9���֜0@�� _o�sTI�oe����bI���/a�y�}t�E��=��}K�l�v�Y&���A�cZmz���B	�`!��Jp[���cl���C~� �<[X�M�TEHk�_g� 9����}����ůCAN��kAN���jyp"��\+q�Þ'�,c&��N��ޱ�����x���`,ˑ3Ɛ�oɾb)�0(��d���Gd	��z��q6��p>�9���eSMV�XY���
�����P8�I�$ta#i�h