XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���V�l�F�8�4&kW��)�[]��p���e���`f#:GOw�����ۏ�Φ[��X]ˀ�j�<��K͖JR���]��E_-ȼ����Qׁ~-���z�?�JH4�!|��A���>`�Xm���U���x�_�J���E���b��8��YT��x�A������A�+�����b�Ro�%��'�����2�*���bc�M��twFxrlˋ����l��n!�{��
9�����P���a|��uF�Jf%���^C����4�,;r��{%�t"U�8�����7��x�7�&q/�<��{]s�*��b�FԖ�51�'|�����]�
��2���[�y vV���a�7P�{Ã��ٛg�������׎!��]�+ �%�R��E{� �V�9�j�ԕ鬜K�`�D���f0�v5��`^��;�r�Jc�#W�єn��v���a�˜i���.�7�?pYg���J���V�uS#�,�D���ny��O�Mՙpڶ!K���~{](�V�@���6�}�QJ!�	t-�z���D��z/n(IY͐��"��pإ�NC���ѵN<691.I6���"��<������#Ȏx�-Uʯ}�Z!����<?{0�+v}ę�Z�#*9�~��m��ZFRUM�[�#�NDۗ=�e����Y>��d#e�]^g���`̤����\�ǹV҂�H���,�*Y&�q�Iw���^�I�Iz ���$1f���5a�9���U2u�=L^~!XlxVHYEB    19c6     900�7U���s;����	���Z��F�9Ӌ1|��w���12H���S񽙺fm�hca�(�o��|��6U}�&��A$��ɳ!}��n�w�� �:��۝��XlO���dP�ͅ�El��k�V�Q9�r�'"��ʉx!��dY%�Eb
[��ɺ>
⣗�j0^U/�8�y3٬t<��H�ӽ���� �k#?�r(�t���unaTi����0�R�ly��ԋ>5��Ecʻ���5O��(\�w)�8������X��ɦ� � ΗB���.��ȧ��"�qң�&�����5��苮3���V\;�%�!'���0!ά���g��)�?A��
D����NO��1u$�I:�k�����Z��t�.⺙����!Sv�Z:�j-�8���@hB��Q䠄����\R��U�}�I1���=�d��n��!�	ߩ�Ku�t)�q��ТX�	��c��J%y��JB��>���X����Z<L0O�&(�w�^�ZFiLH��DTf��p
v
��;�~��'b�^���L���ʯ�Pogf�N��k�m�]��<9�;:�TX_潡�B���>�ɠiRFd�YùƟ����;����.H���\W zf)�C�/����6
��Աj�79n|�4)�����:2>��;7�zb�.FLg���3�[�����[�0�;�C���3hD����C���<���xH,��-���cqǯ��\����(I���N[����J
�E{H �ʔ���z�X/)#�S�[���x��*ex�|qzz==�m��2i>�)۶R�l��\�͜���� Ԣ#@���;��C������/�۔����9�7Bro�6:=J
%҂;P��,<��eȩ�^ƷO%�7@k��-:M����.��r�7F[~G5��bތ�zz绕�#��K��P�T��l�]�U� )�c���r�c���J��Ұw��Ҭe�|���j��!�G_Njw�/����x���ޕp���+����Δ���̢BY5�l ��	Nv$*{\ɤoo�N��-ڴ�3�)��p9��R�d�Pm���6�?��d�@}�,{j��ʼ�\���?T�D9�z�;�u����
�;�O�,{ݣ��y�k�T����-�.�ʌMGɲ7y�{���/vTȫ@O�>�~-�J���s�Xm������M��	RgKx�;ͽ�.�$?�U�y_Z����^���~�s,�"X�_Z�͉oV��ۅo��)���������Z�E״hI,)����'B���E/�	�y��d}f0̆J.��Yu�G�~j�˧�4x���C���?�rl�#���� ވb`�_�V�n��f�Һ��up�*��2�3"��ʈ{��t�Z��Ȥ���&�bL���0��J��e^���������J����%�o41:?�!���0Q�`.d�T!���5�H������!n�ٖW.?�9����K�������y	�u���V��/�<ϐ��_o�"�cs+���9�r�=]ekn�0R���OҠ��6u��&��a��of�O�f�1T��jp�T�c.ě��H���dz	B��ϴd/j�."�r�g.��|���D	($�jAPT�Rt@��\�(�;&P��|S��I��{�	P��i`����%o�"$�Ֆ�
r�����F (8�vH�bV�*������ƯBɓ��.޽���^�-��)q jň������
�I6����=�摂0�?rc����Ж+
����,/7T:v5_oq"�7Qip�27>��m,4t�~ޱ�J��Ϛ�8?�b���\�4Z�蔅���%�q2�S=['>V;2?b��f�Aʄ(�n,�4`�z�A��9�v�t�X�@�s��ۖ�T��Z5�PA'�� a6�{:��I����] ��Dl��n�4��:U'�v^uU�ݙ�p�5�)��q��T�[���F�d���hϫp6�9S���)�ǩQ�783&mJs�9oԘ7�$�-�OK�:k�>@Eq�u����������o�,��}7IE�m+���_�%�Ū�᫤fB<�,n��+B�X�N��=�l��vX��c~�=ɏ�L#	2�{@<��_]���vp��-��O�$��� G��fj|�rb�]_�$!;���W쓕�-��J�7%��gK����J��4Cia���`�c����p&�ýh��������'b���$�mD����n�%DO���Rʡ�Y(*:���g.�M�>\��+�'H����7%ߢ��N& ��4�Ϟv���{���iqw �