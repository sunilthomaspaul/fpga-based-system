XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��R���wf(b��?��n�F��3��������~����^����!�"�r`$Lfc
\�B���:�ˎ@�#Z����n��ɴ^��qxbpa��$9�PG:�k\bӈ�&U��US�k0�C�F":#h�b��m��PP�j���.I�5��4׼!��Ȕ�ų�[��ʘ�$����W7����%�������I�����ᩭ} Ŀ?����+&|����%P������ѡ�C8��
s0$��"C���<,��@݄��I�8w�.jO�Ka*�8�ѧE`T՗;�}v.�c�O4j���]C�J�B�&�>3et��+��@d䧘`/wѬ�kl�ۂ/�����ۿ�<7CBҴZ�c�P���>�����n��Y�It�C�|Ā��$S�|�,~�cd�6D�%�C-�'����8'��Z�p�b�
����|���"���Sii�"4�0��^	*D��w�0;��'�܇�L��������=���f�0������>���<Ӡe�� +�5��E����ȲS���&7�/����4%��[g�
�آ� ;�X�������X�Bۂ�n������[Zi����v���7�z��&�gɍu�UP=�>�;�7;�����@�GE{ސ.<�PS���>,	�ئ�Ώp� ��RA&+�t�lC��1dG'�t�!*���&� g��CGu�-Ld�4K��V���3X�����}���`��դȲŧ�IJ��"f�9^�<R�Ǧ�n��֜/�b�zT�WKm�GGXlxVHYEB    fa00    2620��%���/���~�񾘺(��{=��0�BK����^C�v�_owA���b��Z��݌���*�͙f��<߻���=ot@�4��g6�_�����<?��N����K!����!^Q���s04�k��L厪7L��ۈ�o �����e���n��E�7�s�X@��9֔*�w�Ӝ�m�j{ｈ#x�C��EҢㆽm�� ����I㟹�V�q1����O~yo�A��tT,�=���34~�D�'��Hq��`=Y����y}/Ӄ�g�Tuءm��Wg�������f�Û��<2 ��I�-����aޜ��[3��}��IK	��GcPI�U&���!�.���6B�ϼm�2(.�  s�|ugyx�����H|������ֆH�M�d7U?�
�t�wK���)̎��Z��_����r���T@��I�-s�[?�o���^K�8�ŲHP)��j��^��X�f:	%Ɂ��v(ܹ��`W��~�G>7c��J�K����L�FE�zn?<b@l�s!mǧQ����p��-pW��ݦ#	�� �<-C6�v�U��5��E�+
���Z���Ӳ2��a$eR��R�\s�a��U�t���Ӊ{R�1Ԥ�/�p=��ͬ�H�^R�S�h��u�iy�ٻK@"�Er���m>��kA�W�J��
osm"�_�g\�{h�F����NgE��&r��A��i�x����w��� �d�uu���[e����-@4�z�$�8���YEWb�Tgz{�]r�Q��68���VLO��.��F�n�W`DJȕthw��ʙ5��xk��k���7A����u�,͂�X�>�/�9����e��T�E�77v,1m��h�z�e�Yv�#�<~�����k�Z"���W��%�ng<����8üV��T��G�)�b�V&���ʉ�����*�O�i����: �7����dW�_�j��D�4P}u�B��_�(�{�U-�U�
�e|ccX�Ɣ�p����7�uڷz��\�jX+A��\��e@s��m0�5"�jt�=#��>Z�Y(R��n��i���&N�ˢ	�ж=���N"Y%�IO��9e���9Ք�Y6>kɞ��u;MUr��]�/�+Uy��5�@�#%l��� ���U���<9N�=_���,
"_�3Ѥx�a��̿�n�z37y�(��*_���qW?��(䃕�ڋf@JIN
DJ�;������#ڨ���&��ߝ`V���i3m��t���BH��g9�U���)�����J=}���[�p���q�ܶ}�58+��mH9���Ɠ�9��V1���n+�K�W��1���'�C���O�ے���[7�D6Ћ*ވIK��0W���q+���y+���m�%`34���o�ZVI��G�Ӟ�3	����[�8�K�՟��7��A\/7(x�s����j��7��$9u1�7?��l:��	�ہ� >#���_�ۅ��˥�����Az�����/����"!\���P�F���pY�����DY?w� 7%�yȬƦ���L��v�f���?xFN�&��Em_�Z��4���G_�
���yLDgd�yY�is�|��OԽ��q���r]|C���j(=��v�&���7xQ���Ud�6��p�Lk�-���R��y�"Az�9+.���T�O���lT�U�`B&u��O+/.,b+7ǔS��^�)=_���-��j}u�}@hgL��BU�(�D�AZ�=�g�TGL =�I?l� ,'�b�M�������Y��>ܝ�NG4�����=q�����ec��Gϖ1����=��4c��h�.�(���=��i���/�,E�Q���R�Q�a�Y{�F�!ƽV��re�߾�^����%��N_s)����=�+A���{B�����N����K� ���4�Q��p�9A�Ꭹo�jp�f/�Y8E��!f$X�Jm�,�
�ǐ�-G2GшeP5�FC��h�N�w#9�m�bz�-f݌�=<�I?1�����#��8���Ð����6h��ӄ�g�/;n�[�n��D�DG�m�3^��Z1���D��X�2�zWea�[���y@"�8���m�E`����Q1q��gE���U���*��[E0�(�U�uc�yly���*���$ߋM#<��������'�Ax�Q��%���G���\W�=q��u�a�y�h�8-Ĵ� �����fGx]�'��g�z��1��N�4�w��l-"�"
��'�UtO�gt�1���'Rx�9�E����_��Gݍ�g�ee��]�x�;I!����v����B���:��T��}����[Ņ>�r0�Ο|��i#��������vn��~��,�#.��.��o��2���3�Gd�ՊlR�H�|��R���Gf�+�Ͱ��ei���'>{�[ K/�_�1}G��?߹W�Z^!�Y�[��,%|O�/=�Md �s��K)a�Zyy��#}p4���̓�.��Ayp�o������pe��.m�Ä�8&γ���&��J𓿈[b�p���?����k���,�׼�Vx��Y����4������)U�>~@�</���w�&ʪ����,*ރ��~���	��<JM�ק!���z�2͂�C{�39��17@)�G��Z� ,����R#�ek������/�3�ݡ�����y]���xo㯑�;Dg0���b��Zx;_���i&ڗ뇈g1>�^�S'��D^��f*<�`N����\�5�(���j�}[�!�k�x�7@�3
c�O�a�e�gF�/���Z$5���Z�!n�'��;����3F�qP]����9��Wk,V��ya���B,����
eG�����}���ٵw!"�����u��zI� Z>V��Z�k�r���_uF�<�=,0��',���W0�������N���b�Z6Q�粭���$<�Lv�k��(jjP�����]ޛ�7�<�-.X�"d��p$���Ča�Z��,�����(�x~��
��v��Ã�<��qm�=ل],�~�N�c{2%j�w�>�/�W%�� ��#MEu������!i�{��3�X�=0�1|���(�A��cQ���)Mjj�R�]�O�k����d�cbps`��w�J��W�͙Bɚ@8o/�M���ܘϰ Au:+��֠z03v݀P����	��>�ن�5�B}�RȎ��`�"{��
�n�`%��F���?�8�!u`�'\;/ԏ�7��i��T�w�of�����]ñs�W9�����]R���ƪ)C��I�����u�Z~���)b8�������6���8���e)����ZW�S��[���e��w�X'Լ�$��uDC�_y�3�\�����<�&���
�W��3���|��X�,'fai�>�cHbNF�B��Gp6_?~�*��0s�� }]�����ԓ~�Ĵ �H�0N��ή!TC�l.@��.��Čy�mi�S;�a����e��Xb�Q���2X��r�k����r�C�T8�b���=4
��]���p��R"
�1���)�%�b�҇s��hX�
�3�� t�k�W����c��"������8�~�U�n���ȳ��+�:Yj�4~k����b<F��_��.�� ��rW�x��	��zhk���y+͖O�~�E��-8oK�����屏���k�fhG�5��\kb͖�B�O��<~�W{#MVL֝J�D���w��0>�}���mP�_�hd����؝�R���+L���d��N)6~Z��<t��cݫ�񉥢v����ό/K�a�-�pf7�8Fb Ue��U�� "��6,)c�֔�~%��=i�&��V��ƭb�3�^�2%z�2�����ڲ��;�^'�ї�J�Ն%/�x8+h��`�G�> ��Qͨ��H�����Iԋ!�sO�G��Z���xń8Ƥ�,%�{P�M��S��*�XYz䯶�JLk��ԋ�y|2Dy�(��V���9�L�i2/��۹��Cd/���^�@j�	O�x\G����~b%�{Ӭ1Z��u�<��+��B���I��d_��C����!�vAW����MF���H�`qH�����&`�o��#f�\� �t�!�|��X�P/��>��'���YD��Q�����b�DI��8�h�xT�� S&�n�~h����u���(��i����XGX�E��\��y� k���6��-�S����i��2Oy��=Q�Ĳ�<6ӳ�]@�Sn�ӣ���~�ā��/�t���*ZӱƳ�=L�o�0�+F��W��`;C�TP��^�o����V��=����6�b�Y�����_��9�^����|~|�hh�3 SL��a�M��t��7����]�8y�9��r��u�\>d$Ju[��<-��:���f�^��#��ך���d��m�z�d%�&0kB�� ��$�e1�E� �ƃK�:��%%�zA}Dz&.}3`���O�ftt$0������W�Tϲ�tpb�G�|��7fMtdu�woo^i���⑶>-���=�zW�7pr��:C滃�2�~��+�ט,�Laz@�a vx�0	�8��J�a�y�L+�;򂱹�H(�+f���th�=�q���ܛ�-)��1�pa�ݽ�wǢ���b}{9WU�ؘ�m�|y����v�T���H��$ �Yβ�%haŔ�XXKP�@PgY-t��Of��r��ۗ*���=��{%����8����� ~�/�WW�R(gH��i; +IS�&��zzJD*�#�d�����uO��C��@�D�4��"�Is����6X\�/ �d��f���jdnu~YGsTJG��+�5���.�AR�_�/2��KF�0�����}(�Ob��v����H6�lW?�KAFΉ8�:d�,��H�݋�moz�q�-w燫�����v5�[Spl"������r/��-Q.��C:�4y�E����T��3�E�����ϩ��A��trT��gkɻ|�Z��b@q����Ô��>�V�]l�wfO2����ܼO���]����qݓ�Q����{�18�t$x�{��
s���n�� ���8o= ǲ!>��)�+�&?Y�^�0�`�`$<j��ƈ���\fm�q	#����v{'�M�RV��W�q�i��{�f�uѤ���9IC�XH���%��}���C뛈A.Hw��1[zv���55_�вHA1����@���jk���d��;{G�i��6v3��n]�pD��h�9m��~�V�GOM<��D]��B)��a/�	B9�@��F�EKV��|�*�ԅ��W��
(�F�{A��3^+t�B<]V8A8���e��Vo���Il��8f�*� ^ô�!�ZV%~<���?�t��"ꡐ�c��%!�=�a�O�ks�����_%�_�9��Oڡ�	D���		ԅS&5����)\����^�G˭��+��=q��lŻi���K%Ī�>��Q��v���b�[�-�����i��k�^��`���hk�5-m��6$�_v�r������'�P�i �]�F���vFUqB�p�ޝA���`��(n���3��Ρ���jH�Qş�Ɇ����
&4bߝC�!�+�:`(15K'ܤ��-��රq�c�\"g���T�)PJۆ��`�y��/�'��I͜��x�f���#�J���?W��IW3�G�S��Q|ȡ�P�J�+�i$x#0��?k��w�B}/�:m�2����VS�gK� 9A�����S��)u���PI�'��/�	3��̻�_eTn����x�N���Hc����TN9�3*�	&�=���S�`�i!'L���E"���U��hD�Z��N�'�3?�R��0|���4���,��&��A�~�6qu�7|�>^Ml���T���qM�'��Z-.�xT��ވ�Mջ�������ѽ�(���<���!z�̊g��W�
��H��]vl=�Y+���O�A�4Z����c{�����\���J�ͩ����]��QVIH����N���C-c�kG:Q�J��y/�lt��q)��p�^����E>e���ATk\�",��y>��S)���*X8����>L�<��m5�4Q�ޜ��X�Cv�.�q-r̩@Yf�����b g�6�E�|���kpl����A�@��������Y��
�M��}�A�e"�&��H=E�e#���3�8�Q��>���B�5�� \'l�a1���x�b-L+��n���}T����] @V��m��vD���a+B�j���,s�*�b�ؘ����wC

fS���C[.���pǔ��y��`0?
��A3´�AZKH����R�k^��Q�m�UY�(��8�4$���ꈚ�X�s�	*eXA����^0�-�����dS.D:7rH&�.9۾y��H�L�Ĩ�O��Bv^ "���,m�W����S�]2�x��I���������
��7��S�n6w8��H��t����s� �'|��'�8�5�~����+�����>0��7#�5se�h��oӘH�sE!=4�rHrI�S��Wo�d��'��¸hRg:y���9y2m�k��L��֭k�C/��^�1�ۥ�;@�\�B��}x������
�&�8njX�IS(j�1t<UIl>(G��������w鑝j�b$����$a,:�zl��{)+얝������{�E����q\1��F��S6y�n�̴��Ek�\\���L��9R���5%�����`hQ�
��qq��K��`�N@��U�X$J��N�ߛ	��Wλ�R��bM�!ݩʕ�@�Oqi��:���JTU�lɶĶn͂�L��>a�Y�~!�|����_u0��$��HA��hIOk��G\�!^��'i�A�ğr�9k@Q�Q��v���*j�?�"�K�X��n�:�nڞ�j(��%
��*@PI��n.-{����n�]���z�{b9(SK�+ �P�U4�i-նx�ƚ�.n�CcH:�����(�h�4ܞbJ#U�����|��h���q!�+<�����6�a���ʚʼ �|��ТÝ���:{��ޜ)
J|Q� -%�����5f_�����*���g
FBO� >���Z�i��Kr��'��1�i�9,s��FVu"6��H���JX���f�1�St)1A-�HD�|$�P��z�;�.Ӑ�1R+�����$�KB�m���ez��������{6K9d�&[���%\bx���t�ǹ���?�o�%��,[ �cȪ�"���~���f����C��%�h�j�[*�ѫ�v�m��A�����͔�6�����^q�[�(D�+�����TΒܻO���6��
���_ o���w�SR�Ӫ��V h�)\��	b�L!��͑[���B�s��y�ؗܟ��Xb��=2�XA�����OTU�f´XW���5�6;#ynu����铳��u����vRIz�Ha(�Y��̐>y`iy(Y��Hm%�ji`7���[��$�ky��̑��[-�Vm��yE!j�\`�W��)�X-��?�rK��WK{ ��U�"��2_e/a�2�]	�m,*��%L����`� ��?��Yw^Z�)���Ö�@����X#ZD��N�o�T���H�%O���h&*�aE���O؃�Qq�ٹ[���*-���?p��@ѕF�yM�ڊ��h�h�d����T N*d�Q�Ԇ"�b�8�0�u A	��:�q��II�!����Jխ='��j�0ۏ���Af:��]yV��J$S��X�]�T9� ��}0X�r�͒��S�ύ<c���(ET�b�D$?�	����-�Ή�� .�NX��6�J�O?ѷ"$���V�׍S�D��;�Rc.G�������8�������Pϻ~��7|^$�n��ž�C[s��,o���t/_h�k[��H5�U(���
���~�����ILN��� �{4��xȀ��O�w�b��tM:8��y��!��S��P�3~�����4�k [u��3�ٟ�dF6���m�Ҿ{�_6�L2ve�\����z��,����M'�����J;Z��TG�4 B<�����\4]Fz�Y���+�qP�s��7��fBh�o�kԽ�P�Wk��+�|���M�8pp�N��?%�W�⛉ �5��T:�F��V��g��"	�U�T�35gA�J��zL�؋FR�P�|4ץ�4������C�Ք*:.�#�=(*q��� ֈ�V�S�ԛ���S#��C�0�ʢx�Q������ձ͖N2�튔��y����suS��/x�\��l=�1nL)����r[ ����ӈ�{eL7GSXFY���o)h�b����j0��k�h.,���W�'���{,y
��Qtk^'n�Ք>���P�H�*#���y���k�GS���.����r��s��^��}(M��_}���Ȅ��v%���$�Kq�03;f{����U����S���O���,wLd�y�i�ї������&��:�i�c�XV 92ǌ�9�n���@�+i�\�IcZXm�p[)�<s-g�pq@淩�O}�ǎ����n��mZ�b�h	������.��¢J��K.x$	q��n?N��/�nl	�~��D=*� � ?E(���S(�f���񍃨vM�eX-]m5�(�&���Y\�k0��S��=Q-��\���kj��3	�����W�9:���%��X*���nOΐ >��5�O�׸֍w�ށ(�ئ
���B�O_	m��ꔽ��a:�nX���D��!̢��KCeh����� �G�٥� "�p����s�t��څ�jJ��a��^^�Sj7_�f�Q;�z,��׬l�rANN��i�֤�[��C+�x�^c�i����!D'!��6/���JL$�`����/%�����x�3�ҁO���e�&�G�i�4 ���:-�^�e~P�-j�P`�Ԝ������������]n�He5� �����8��6��1�o7!�!��J��w���A�ס��JÇ�<h�oh�Jxp�_>b
�Ɠ�8˴!�y�l;}�9����Z�e4Qs���7"-��>�k-���e�~[by& *N؄/�ꖏm�f^�Hç5�ZE�Ide�E�̰nG`b�Ԝ%w�����E�7�	������&<^q
j�A��W�m�22��a�7� q:����[�PJ��y�n`.������w�~��hb�?����p}�@1@��w�+.b�V�� ���]�׶�|�@��p`�D�(�u�����u�Xj�x���(�Zp�4���\WPO�w���Ϝ�8	��C���߱$�z�Y�Zzn2�"O�����x��[�K�e�: ɬ��Y�߯�p"1�'�@.�|:����~��$u��qf��K�_m3�m�_o٬�:�]�p��*}�Jy�$���*�9	���`���N��f�y'��0ҵj�E�E��JK�#����^�'f"��cp��Pυo���Bɏ�ѫ�������C��7�-�ιJ3'X��YR.�qTA�̎��y�T_�+,�Z��� �G�G��8�	ӷ)h�*��H�:e^ƌ^�'�t:�w�(1�J��/ߑ����T�8ԏ+{����nD<����P)z����9o�bXlxVHYEB    37e0     ba0��Oӛ�mV��`ЉI�"c����Xxv��z��>Cp	_�8RJ>ʲ&�s�G]��gx�j�RJ槯uΊgVҶۻ�o��{Ǝٴ��_ғ&�"^:�S��!�g�:QH`�4�+�#0t>ꗬ|��%6����=T<g��H��!K#��+�m�[�p��f���dVЕu�R7~����:��Ѱs9g��pv�W߇=��C���P�0���нx����E(Q�3#��x�F�H��󓗩e�S-O�xm�����WDɒl|�ϫ}��� <�;�k��5�,����5P�v���֕2k���21�q��|�̬�8,���t:#�߅<*�{c�f/�rx�B��&����(C�����>����OL�%VU�BB�w�+��-KB�U�F����/����|���l����MQ��	ªu���x���˨�]�YIQL���L���G�X�Oc��������d6CZȮy	>���
��Ūyv��(M�P�Lk�5�$�V�+W�Y.W8دB9YoK�N�61.H U�y2�f��di$�V�ؐW%��t.oF�ZN���n���V����3��>��Sf�f U�>�>
��`��F}`�q��x�MN��}�����`�=�D���说(^�H�}lt���<-8?���
rtl���7�Z�;�����Fr۴�(�:�TB�䢘�댵j,�'�>RЖو��+�ڐ���\�MF�O��l5�Fl����ɗǅ��/��Mc�2�h�C���lvB?�Kn�<ID�� �j�"L<f����Ѩ"L�Jݮ��ëʥ���I�h�|c���^�W[�6�z�T� <�ڰw�*�?���[�"��;�cxA��5��?��'V�=�{�5=C�r���8����Mn�Ԁ�lO���\B�	��r�A�{z��6��Ln�+l !g����-$���SRJ�j�>������ײ�3�W%8�}K̮s-9�pQ���3�˽ߺ�܉TG=$�}�ױ��\��*���φ���6.|�!4��2BeA�Cl�`�J�������i�lU��в`v���A��8��NV0C�V��0%�lK�����
BYz
���}��9��!��	�0J*E��+�~R>_r�	D��
ZU���u��E�v�4�(@���z��C�)j�̾�D�A.7�3�&�o|�	WU�+�0V������q��$��Qe��<)����]��Z��$��v��o����ȱ��U_I/4����PX�L!��&S����0[%�ee��U�!�A8xO������|;2��ls,��������Ճ�`��L��k[z�P���$�%�������QX�\S�Q[6��
h�~�2������c����Z�-���Q�M}A��%���\��m�`��Icw��8�.��b�fo�i`���Xޛ�c4L*;3SN�B;�N�3rF�J�¤⎾��0+�b��s�jYH�̡���5�0�+c���ru������
,�I���4p�������m��x���Ȍ�,���w2E�f>���]	=�m&u�%�"���A�a��r/��Wx������ҵ�`ry/6�uwtiF@js�}U��L�{�,I+��[�X��e"�jQ|��?V�
�v�� О���i�$J�rR�ho��H5Z ��f#h��f4L��ݍN�Rz�4hB'�?F�6#z)����Ud{���9:�4E�Y�!�E���*��k�X�9��2��Ī#i�6I��5����ᤵ�� �ɷ|0W�s<�(,���2>C���������+�R3�	�^S/ɦ������A�b�cH���	bMs�ܝ�x���23�}J�"�yB�XZS��hyH%�{>����d�`�BȰ��{c*����!����1�Z�K2惷F��"O*�W�2�B<4v�B\�R�,�T�5꧍nxG)�
<���n�^F�"�e���$@Uq�ӱՙ2Se4��FU��nq���aZH�Kv��� ��A_Ƞ�Sz��������#�f!z4Yư������5M��F�+b��\gW�Qa(�Xok�<
�	�+3���-/��U�f8�Da��>4 � ���Zx uI�kg��1�Qף��w�C!���L3�X�^Kf�%�<B�]����)�_��Lɸ�)��j^�B �X���0���L=@.�p�O{�<D}���n/��.)j�PO�i[a�������}C���p�xL�DO�[S� �2����j��G�)�ď�R�R�V8���O�m����ĸ#��hY�����"�'z~r�,��E��UoVI3�P��C����m�'�i���~�W�G{b�<�mk�L˚�{BT>�S��0�Ī��4s)$�U���t���+�~>�Rw��3�"l� �Lme�~�i=�$k�f��?��Pᡈ �:'!`�.�on�@��J|�:��7�iM��'~S�(�
t�r8K�6�D�;gKjS�R\\^~V @�'�Q�l|���||R `[�֊����sVd�u(�UB�{��聛@�����m��7|p�֡!�7.=\h�qY�~����n-WX�`-��f�yo����*�cP�W��:�+�%����U^���7׷�M�����PT#���7�J�X������Æ�`�^ކ��Ccѕ)$�*?���X`p�ȩL�pZ��W�~5��Qs�aa+��y�x6�%w���Rvы�w��Xk�9u��l�u~������;����5[�z� y�w�c�aJ�`���O1�T��;-Sf5�yL.�"�=��W����N>�Nn)�K�@�����7lu ?���D� (,S��c�~MVf�ʦົ���
4n����Q4a��C�K��z�vv0jT�<�N$x�U�֝n5 ��e�PH�����wj�v)��1