XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��=r� �ݒ�[��(�L�u=TE�3����ɀZ�":?��Pvɐ�W`Hg��I}̽n����^Tz�>ߙ>�A���ܻ�Y�'H�G��b�W�Zw�"Z�
%n�/Y����b��6=&�0xU �B�#jU��9�{�(Jn�6������U;ԧR�Iڽ���`)}����w�m��[lq����T\s
)�H�(4H'ŧ��m􃇦p�[���>v5�9�i�m�7��,=6擧�V�����yAA� xұ�����ߴ�~��m��:49Iv��-b�,j�2�w��@[";>T!���(��!w�2�nݕ����~LU,a��v}��"��֔��`
P�ޝUW&�e�.�O�`�JIZ�#��|'�n�����ӟ������P־�_����.K=S��Y'F x_2�?�Q�{���*���
��w+�?��*9�n{��tB�덬;T[n���P
��o�f!}�L&�qe�.nH��:�6b�E��Ø�X�O�4�MO!�4� �*�\�?���Z@�p5Yrq1���)b*����I��?��G	��\��o}B�F@��{ӋPf@v��"�t�(
��k��g�5X��G]�kgZ��g�CvF�f��)>sl'�Z>"i�G�H�*�TH��t v�Eb�'J���".o��,����w�ڈp`q�ooG�g�1~��J7�KҫWlӔOX�t4�8F��~4mxB}�dw��h_�u �����)�7T)ƀ�)�'��i�/�}I��
�XlxVHYEB    5571    1410���:2/�c�yzo#Mqi���"�!a/�V[�B��Y�Ɛ�M+���/� ZS��XL԰+SӼ�_���F��1@DPxD����/"�-��Xg#5�����z���Y�X�������z#Уb �+@:��ԛ����.WҘN�G�	��(���D��Pp���ѕ*���Z��є�De��aO>�c�̋�An�!���)�Z��1�V=Ck~`�l�k,˔�NR�J�K�~]���w�V;D��7oV-���T���I�e0Fp�����?���?d8	A��\�Q��Y��A)�d��ts�6��{�C	��D��G"%[�:�P��tC��(����NJa��e#N�>aX6���u�@3�?�T�򫏮�rE�"�1�Z��*#٦:�fj��@�%Ԟ`�W)��0/J�k��}SFb��\��|�	B�9/�~y����5�~9h���֨@���z�q��d�UP�2��Z����ɦ�2�����^b:с)��?��H3b���EK�����/��'��d�ꥵF�i��Z�)k�E�L�{[o���G	�����Jl����ed9���13��!�
���`	����,����^$x�1�*>�.n6��;��(��i�͘��}�xB�$_�I�� ����N��h���D�	0���M���s���� S�/E�ȗ'm���Z:�&��{�|6�2�Xô���!8Qưt>�}B�����d�|;^n~ϰ��!7
�}�{
�>=�5���������i=��B�JN��+�*��)�(ͣN��s��y]�XS���PQF�+8�cM��w\���!v7}Ԅ�B��L�RY�l���������Z��~��@�|=���	�P1�b���nϷ�@��\SN"q��ԡu3s�Ft~����l�qJ��!s�-5��B�~sf�Ǆ�,	V�ć�%8�RM�'ھ�o���H�5nvà�RVh�����r�ۀb����%�W��gZR�o�l�i�OM G�J����8!�2yxg������Eo7�h�53ە\#�C��ڬX��0M�`�a�T�t���?)@}�n�Cᷴ;FkI��J������ͥ�b��oE�ױۜ��"�Z�5�7q���@��cY��᳢B����BMG(�D� ="����"�!ZJ�K�Ŝ������B,A��U�phHJ�4���sI�&�jD0K��↊
֙b���K��u�<RO����5l�5��1���e]cF�������Kb4�&�����%a)�T�����$�aB�RVd�^���LMb?��H<BU���r �R��������*ⴥ�� 3�|��9�>��'p�yV ?��~L�l�ܒ�O2��@����E�;�;�$����4ƣ]z��w	�Rߐ�M8C�!ǝ}K3���z����ҲQ(������[�:�,u��e�d7e�ΪN�����j�C���Z�����	�k2��	-���prm���Ng�w��c���Z�7K.�F�+L����%������my�`<�d�5�d��0�3{fm�!@?N&���.�4c"��M������9���ܘ�43T�0���{�#������SU�^����kj7N~�~�Ԣ�4R���P�І)=d!��ۊ�R�;W���lT�t}4
I���lWtdNPhol�yI�/�@�6[�|����I4��0+]�U$�] �����eTG������S�4Wuܿ��q�w����=�l���mɷ\�M0�����=㶳��- �j!�a�Ԩ�|��+݅��ui��������<�[RE���Pt�k�����XKpV�1�B�pSƑ�g���[䎱j�(Y��]�ez��~T��J>D��u���?�H����V>tj1р�MLP�PG*B��5���`VZ���*���>/���}�C��?zb���x�V��{c3��f'J���>h����u�S"J��FG?�?[�޾p\GQ�𲓳3�B��]-��ٛ�o�m}�zXZ/�ؚ��:>8�,�*�OF�D��ֿ��5��=����e�O>ؓ�3�T��BBy4#F�D�>
�iv���;<�D��Ȁi#��;n�-�vN�g��ο�*�Zi��9��n+�SJϠ�O� ��� �L���.+7��R�t!��y��kJ�%IDS���rͮ���ᩎ
I�uFK�
�������>{G���Y�Q�oA;�����@�j�F7��X����1"���/�A��)�$���7����L�Q&0T��(��;�*j�-��ң�j�0U��Kf���:�β	=��yx����Ѓ����ВQtt��xnz����7�I����1��I�5U��4=��Qgq갲�C?��2y�4b�W�%�&� ����C��Ln(q����4�#;]ojR�V8RJMK7��?��4KF	��bwCؕ �2R�ȧ���J!�n���N>�๫��Y:Q)Ԁ�l }��Hko�|>Z+�:��S���6���G��y�6���q9��s��2��3��-N�5�Lh���ʯ��^��3ȗ��]�� l��G���H�$RPc��7?��6��ڠe���\B�k�����*w�c
��y�FGR,X��,/^B�k�'������pAA��*���C�'�~�6@�e���v�m���"U{��B~��`�s��=Ų�%�,B8�r�C
\�S�JM�
"���;��e��I7߇Ab�;�o�Hò2����A`�%��ɛ̆!M�4ѝj |�wK�j�'�H���gIF�>3a��u!LKT9�j���ܮ�)L ̩ڏDƋn>v�}h?)7�0X���*v����5,��Zs�*!�-΅�}�˖�k�u��u���p��n���1�c���vu�J�ʀ�-�H��}�'�sR��I�e�)6b-CUZ�`��v^����"Q�s�	@6�ţ�B�尼a.ƭ�R��x4�tE���y��Jj��J[#)���#0�ԏ��I����_���UF��'o�Ž4ʃ��)g/�����+G�Г�����`j���ÍvvL�ʕSZ_6�mιў5��e)�e ����ȡ%*��$M_��9n$=�J���P��BA�7&J�>�S��V��P�tV{�Hyp��m*��p*�t{Df����ɑ��н�)щ��ro����G ��6\|W�ͥ�Q�HKȹ��iX����zsU����;T��ʛi���_�°��q�R`	�8�(}�Ǆ�ٺ�Y�,���|��/�jҜ�3W_pY8�0���#��鑃���PT�bQf ��,�s��׫	ƕ�H��]2bwp�X��vg|oX"
�P%��(����Cs�Rf1$�<=ր�/v9
c�.�D\Vd���R�?S��4�W�I�k��&�b	�V� ��lܟ]ޔ5yc�	��+�=,�5h�A�r����d������=�{g���Z������s��	Fժڋ���9�t����&k��4<-C�6��j�W����$(�gx���L��n Ľ�a����4@�h/�b_�5�u�����z?��@J�]�����M�8�G�W�V�2�B�����Ql��+C&�������U��p��@w�����
���׿�5��E�Y�MDY�5���+�P��}y-�=��%I`�Q�a�t���F�9�
�IJ��"M)]S��>򕇪�l.�yW�^b��LH	t�����;�Jt~h:�R��Ah���H>�`"1��달��-%�Y�*�3�F�7�P~'&�L_o��i^e�>���w�jږD[���qR��W�ⴍ�������|{Ma76���QQj\�k��k&�>�����da��m���5���K�"�B�O�����<�B��� /c�(_{{r\�4��1��äc�&��g��E����r������ẵ�&A�$�2�o�#4��&v0	����1;�2��:f�}�z���^�h��
����z!Y��ȅ�����D4j�Q"-�wy7ذ.�*��|a9����3Y�)�f+x~�|C�������:�os硰�"�e7�[��.S����S����p��w�@5z*ڱ�ʻ"�f������Īڗ�g�[ �?�,�i�Q��������fI n��i3�"|��!�z�ހg���Ϣ�3y�x
ѧ6?�;S��q��:xA�j��F<�M�ﶸ�s�C-�٢TD�]v��DWBh�Y'�@vŞ�����'8�k�7Zu"��Ys}YG�J]�u�8�R�~*%@E�!/��I�3�^��v��k��������AG��K����;4�\ַ�hL�3x�ؾI[5^����e�0?z.�9���3!
b�f�<�]/�4e���3`3	���F��:nU1Dy��o3<=DC��s�;T���\ �_aĝҔ�d �i�z�4��#�1�y��d�v��TA�{�ۣ�a5�%�3�����:9��i��v�ۿ)�e���Z��{����l̵����j�Ƃ�6�zca~�g[L�,)<�[��<H{�J<0K��͔�7kK�m��O�����wHهlp��U�\�A����$�=���qW<8�j5���-����M��J#�w�Zr���_D�\#���n�ʾ˪'�J��I�\,�]��YUk�T|�p��I���>�ܰ��DW�T�4S>8��{�|c�LO1Q��-���%@k=�0�$���C��&(�����q.H])�8@�rԡ���z�Z��Thӑu��sDsް�1|5=ө��-lqZ�q5�} ��)Z!p��P�6�/����j
*�V�*��8"�U<�>� �3`++%���'i��d�RӼ�e�a�#y����TMDa�b�Lkt���5�_�NI��h���&� gH��5�������U�'�1+oI)���9���e�6��o�CE.#��^�x8���ِ�Js:(cOvm?ZzT�;W{ްs�Q*�:��YF�UW�������R��Tx>.
Hto m$�nቭ8(��䤼��d�����6� 6��p��"K>7����L<M