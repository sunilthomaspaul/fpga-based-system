XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��;a�oQU�$��2$�,�,Z�h��&"nƸ�C�L����{u�r����ְ�⚻��;퓼���C,ն;�Z���k�*��i��3;~�e��>�C�Nu�9��Q����9%����p�؆�"�ф_������{̖�x��y�S�{�(�y�B� �D'��)�M����v�f7Y٫7z&�֜�ǯ��5�������Z��(�$��C1��]���|�.������GsA�BV�sʬ��_��9��K�@��<��F����%wػH�ok��jH�LϏ���?A��b��r��82t�s�ղ�5���]Q��
0h��J�_8$�Rva)#�nWk����{��0���Q���b�o�:>C˷2�/mכR�t*w��t�}rv�z���+f���T�x��<�Ǡ��ؠX�7*POL">J03�W����6�	�m��y^i��~��?�
zK�"Ċf�����&G�Dd�6k���de��d�l>h�%]Z*�k~����T�w�$��#��OzJ��L�M:�%��?�w����>h@#�ʍV~����Nr�&�(�EG�Y$�Ŭ`���� ��|��#��d>^+��0�<s%Kȱ����?S̵đ���0.C���!e9���l����藔C��r~�j�9or������l��t#OC��Փw��:�c�(�`��J��{h� w[v|9v��w��V�/��8�L �ot�	s>���x�������lG���\��CKh�p���s�nXlxVHYEB    1854     8a0�P�׃OW���~��>BY���υG�w{�<���Q��Z�>5��s��KZ��a�L����g�^�J]?�W�a�"��G���[�2�4���ى�{��5�[:�L�xk`��5�b��b�+H�	;�n.��^��^��H�a�i�4i>:YI���4~�%�q��g��W��?ѻ6(D;���)���ߺ9�.�܆���B$OE�3>�P0|��֫4{�@�V��S�j�O�и�I��(.3NQ>�&I���u�͉�r�U<��YB�z
?�[��hW^H<�AE{i�-!�v��*a�`�+��I^iF�}�j�z�	x�O�)6���d)��X1!%xX�^��K�vh��
�����91o����]�f��/ô�B=|��棑�1��0�ir��E֗k8/p�9���Z�
��>w*�zb;�Ȋ~�Q�1�uړ%�s���U��_����[�WD.b�N���P�����%�t9\��u6�(m`;�1E:���[�,�������<�Z�p��Ta��lX��'f�0��P��I�?�f�y�i$0���#?t?�	�`�-Ha�t�=�����n�C�[�Kq�8Hܭ%���}��h]��!����i�R�l�_�R��]�=�A��E)���%" ��V�)���z�5�?�r������'��
�V��e̖�of��?�=u�ʹ�ʞ߆!X�
H@Y��u��mO���)�G8y���<%_�q��&Y�����������c"�rV�D����Z�&�X�t-x�]�zPΝ��jc"�`��ȅ]�Ƶ���d׼g7�܁���.��０��2O\!m����{�ɇ�)�۪N�@T�[������A��b��7���ʒ�qnE9�3�e��K�����^����jsi|�EA�(�a�F��&p���ϰ�#I��Y�a��W�6AJW��#����4}��} �/�:<y������hj{�[�~�+yQ�M=�/��R�r ����˥ߡ}��͘���#��N.(��l����Y	g�ɓ&�Ј�����U��"��_��.E�o
��V)掖��\�����FqH�no&�
�W�pw�2�$�+V�(}����1`k�:zO���ݣ-\SǷ���/����p&�cU�-�?';�Dps�M���A�s��mp�a$�{��E�����NP$g��	G�ל5x���!����xΏڂ�C���n �/�Yb����n�*��\���ti�v/>���^�<��X%��ʍ鑄'��e^�2��S�g��v5eHi��91:n-��^�D¨{���9��Q;X���b&Ó��J��*C�� pJH�#��x�ݒ���@�ZV�-���~]܎*S����W���վP�*F5�\2U���I�s��y��C����g(��"\���/�gT6dN�ϙ7|��)��U�';_�؃��~�ks�E�q_�0��#.ݹ3!z	L�b���JU!s>[#���>�&z�D����Lg�og}~F�+cֱ�=�����^��Q ��W
UM5����V�5PL�Z��2I9��{9(�+S�X�EbR�#�L�)�m-��Ytm}pA�% ����	?��i^轏�~���Ť�d��5y���C}��׭猹PbQ��wJ
^05�w�o٤ȼd���R�B�ܠ|ۿ?�̧�������1RL	��+l���?P`�s�1e{)�����( �#�����}`f����R�כ1�@3E�}�5X�c�
�i}�|�����SmޠWM0Rُ:��Lc��4��X����z>Ǖ_/ ��B˫�h��8�g6	��ٽ�ڧ�-F$է�,m�4�J��ӂ0�^˺�nY��yA�I��]�Q^���I�mlK�+c��\���X����Qߖ���)�c�/Í��v��g6��*�0x�2��C_,Z�؀�p]Бj���C� Xz@_|�L�(ݶ�e?���r���#�h{߭y�c� ����6��/"�4�B�~�]�#��G♬Ԕ}&�h�Vj�HEpP���r�u�#���ƚ9]�4N��2Oz��5����Fn@���IE�qeȂ�j�>�`稏�.�h^R\E��4w�EA��=��kat�6~Z(IA�٢�	A�$��{FLs��|^99��M�V� �ܥ!iP�^'��Dws��$i2�FqjF��7�^w=�}^K�o�J�"�$irT9�C�