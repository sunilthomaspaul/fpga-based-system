XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���Sd+�}��%�4��&�]e���[J@�v�/�n��F���Ն��Ρfx��Pp����!�: ��K\ԑ[���԰�3u�M��=|����@#E��z�߅��5�9��%�mswS]��ez?��3�/zȋ;X�e$����Q5g�(������g�
�<�6%��(�f4�t��>្�Oz�����_��-AZݿQ�[U��NMGɒ��Y��<��3iR�.*����L����y8!JR��?;�e��̗4v����Y���UYdzN,��Oі�k�s��^^3Ph1��Ǌ52�Y	��oX�0oP����c[b �JVg�胎��	
������΄����f�z�l���]����C������Q�+K}2�_��2�$z��V
p���]������m���x<|�~\ĭ����]��QC����o�t}���~΄���jZf2ܺ�:B<S&,�{4��?�*�B�W��D$�(n������u��H��-�o�ղn��SOyѠ��&K���.6Ngqt�/�8А��fC�8I�K��a���2���3��I%��E=�u)v�W�_b�aEt�W��K�$Vl��~�N`S�t�D�!�:g�<Q�}C�� W��wŃ?I�V.â�&�ʍ��6$=\�Z�6KD��=s=A�Y��ElF��c?���~���x	��d�<k�,�"�Mi�=+(��B�jW�+��㈬ ?ݼ������ݰ�!�����I3&�V�� TYZ+� _X���I�����DXlxVHYEB    1111     710*�>�)b��DŲ���@G����!V��V &����� Y,�M�5;����q�T�P⌯�!���J}}�7��@���bk"�`�$sd��e>焾tQ�'�����(�0o��ŉ���n=�ެ�O�K֠�Y��qVA��t��˪3
XJ��21)x�L�ݮF�E~�b����$�G
���۹WS�DH�R�}ǂӕ{�a @����$����v�B������wGJ($��ipQ��$$�U���	�/v�6��fj�l圢ڌ#�Y�O���>���
G�O{�HD���2P��T�l��K�dL��,D;׀>�˦��=�vM] ��FD7�p�P`o'�u������I���{SŌ��L'B����E	sI�Q�U/�䦌��q�ڿ�x5�1:���^=Κ�m�Q]C|M���t��@�v��A�w�	�D��=K��i������"9T6�B7h�u���Tr�E������}S�\��������3�%��M�����ڍ�)�D�:l�+=�B��������/q�-jۖ���j`��7?M�P�7�B�Z;v	uC���[%��E��/�o8��,�V\޽j*<�ӹt���3LdQFm2b��,�;T���c,�6+&{�4���l�F��>�<+F���8�ug��0�����(���'&����F!A&q��*w/^� N�`'���ʑa����Ykw>���2):aF.�{^~�u�P@�;�cK=Q0%Ccr!lC�����n�4Yi��"�Lg��md8(R���<K_��Z�z������.	*�'� �@�W����5�r�@܆Wo�:s�;>׀{+n����DBeo�pn����.�ZW�N28kX���M�l0^)��%��?��g��(��.�ܡ340|��~��}E��3 ��|RG@�$��h�����5bX�ʧu�Ɋْ�<7�Dܤ�gW�q�ֆ��ih��c_�*��\�j�}�z�oe�B��~A�	>H�|�]�gv���u��޶�.��D�+�Zc� �aL���3��qv}��c�l��{���� ~k 9S>��M���[,"�LX�D��p+q�iD_8"�#ʥB��L�"[�x"�t�'ME�p�޷Z�iE���_�!*MD~Z7�ɦ��ek����
mJ]?u�/fΦVL�5���(�c'ן��P���_"��s�N�ʦ���5vv,()���iL�2�|�����_�ϐ����T�t�2��<3|p�~��݇��rx<b1�O���{��β�v�������$��3k���E��%F�5 &]�}�EiĵⰗh�{��m.�^ ��D��Q�ԫ7�pL�j�~�q>�X��a�Qj�e�˦ i�q�b����W�Q�RH-V
�_�{����-��E�����ڳ>V �i䴛�\mL�-����ɟi�2��)+�9�Ɠѓ-Xq"�*������hDHT�FvN�]�T��<�z�M�Z��u��;9`���?���JT���7Nrc�7o���s�	��l�%J�G8�b���	k?�� ��=�V��ㅅ�ςR䔙XMX{\�3��f>:u�ɋ�[�H6�1t��E��R�
�}r�i%���T��O><r ;K>j
��y#VC̗�%̭m�<a��#�w"�) 3P�3
�<��Ҹ!r*�3�Ē��`�ȉ��4£�Q.��VT�b��L��-�E��8����9i�G����N�mc��$�c��� :g��Ԗ"Hm�L��@0�r�Lxƺ��Q5!��mW��d����R����}��~��z��-��q�I��y