XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����#p�OC�����7k�/�t`����	A�8ʧP����	&��94ll��%Y4��1��w^ְB���[t�KP@�P*{�`&a�x���x�PQ��Y%��M�zw��-��4��Ƭ�0F�2_�u-��ER��������s����Zmt���R9����c�֟���_]�J��D&~�a�>�ɵa���
5􁖨���r��}��Z�Y���s�%}�Dc�6�̎���t[1L�J�caqDhT�˫C���9��������g�������x i��=L����֫}��x���ow!�{�oz7���3m<"5?଴@�XRt�yE>r��r^�~�f�J���8`�A������v{@�p8�-G��l�m����ЀK��^^��:��Cl�\żhkΖM�X�7����YLx���kR�@3�9l�aNѬ	����R�5��p������M��[>PL(ԊD=�����x�H��{�;�.}���Y�VE��چ������-\* �V�
+�l`��.�JI��^1�-�"[��"�$��OgxGZ��]�&��$nq*�Y��r�j��0�zf�JP*P�/.MfgSa��4�-us��Ќ8�nJ�����n�*��5^4]��{kRo�q'E���%�&�86���'ch%��&��P�0�
:�*�7y�PO}��f���k�������G>T$'��IE���D�j�ʷM�R�\��5S�a)Г���}�S[ �Q�f��BxXlxVHYEB    1854     8a0׬��y��vK(�|QײX�X�"IK`/��D���R7ޡ��:�!����ái}��ާH͆wP�I�e�QV�Nx1��/G�˽�"�2��Rgfj�b޲������D���҂�:TB�BԴ�� �`��=�m�戬6��;��$*��x]�X��H�$3����;uQ���n2��;�4t���V�!���Kl�+����p@gt��5:[&���E4h�!�@;%t�P�u�"���a3�O�� l�pO�K��`8K�l��8U"KP*���ܞGz��Mx�_�;����Jk���益��.��x	Ͱۨ}p�*�D�~�����B�VB$|}l��m=�̬.Rq'�F���	)J�C �E�hFq�ܦ�ZA9|~ʡ 1���o��G�Gq��H�fm~n	�AT��AyU�b ���j��~�#vf������%V�n_���5����_�x�at}C�W
cg�1�H�]�c��ܛ�7�qI��W�\�0��@t#'���9���	�Ram���e�=F��a�%r�)��+�p��5������#�S2�6&z�a�'��3愌�4nwc�d�o�{'�a����e��T�_H�R�͍o�PX�\�l*���%�b_��=�dҵ�V�Id��k���3��ŏ��ϝ����;���\5�:o1���󡭫>'�l��틶L�an�3��Yp�g�?M�QM�L&�#Kc2ġ�ʼ!�tf�ٸzƴ���������ٕ&Q�)�te*c��a'�6�:)��2�"��z��A5�p� s�^0{֒ʳ;��c 1��m�&9��5��P����Ƽ'�ꢄ����U |V�?I��M�	$��J��%�6����J~�MTF]�M����=��>�=��@���!���)��O־���0����<�7�e:"�������O|�շ���b�$f�}�(�!�b�hN�0�)�Q	�g��
�O���r���G�k��	��3'ƨV��-�p�х�v�TH�������d���vY��4y�`����� ����ϱHk:i����a��H��&ri��~��ܟ�ex�MGYi�W�r"|��r?x�����c�q�잃D�M4��	MI��-��/�<t�-2ˎֻQ,a�m�쏽c��U6�n�y��`UL�zqO�G8���k�O1�ߗ�Sj~*.�5-fg�����n������@:X�p��A���Ք������F;Аz�O1��P/�[����Bl�c�c�e�bG{e���� "�T��6���A�B\9�����u����g+�M'�;N��J*��k|w��ۅ�����D]d�s\�Q�/�:��t����惡�=�Q���R�E}ר��b�5���xo-�q����`�?N}]^O��q��?^[��=�s�#yNh��b����+�@�V�^�x[؊�Hݽe�ۭ�$�؁�����\7�;^DJ=��x2�@���'��:��(q</�����agK&�ز���y��ɖ����X�XieHW9�I�a�b����5�Ld?^f���J"�>�Y��65�}Qb���۽.j��:�ՙ(�_�M$1{�gk�	��%ԻAv�_�N>r����¡�:�)�Q�P��5���Sa'�C��t�ܵ6�&VL�xw�h����Ʒ�1L�����"�s�`���Q��E��+/}G#4�tm[8��R�k�����b���N��N�г����9�]z���T-���Y묌��بh�V�Da�m���`�KWt`����H��LTCI��c���8"�
�)��-V�������&�	Eq�~��ʹ�)��������R>���MǦH��C��Z�/�.�T%�J��G���%��p}�˓�12�J[�`�砘n��g��kR���	D����A����?�m�g��1�ht���9-O�q��Q��O�?����bΝu^��l��G;��kx���t|e�Q"��T¶�b�8U���gi_�v��)P�/���)�I6H��x�PE�nOY?��-��M"{��J�L1�aG��Mb�z�ɄK�\L���A�ڌ����&I�������čf,L��ω`$%A��xuH�.�����?L����9G�M�AX̊"����mK��&��t��^�AX>��G�0�I��L�_͗k����