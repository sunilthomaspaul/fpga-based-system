XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����v;,L��6��ؙ8h�DH�QBY�dp<d��@�{��{��C��O�M�
�dti�Ի6��Yy6!%�~��~Յ��a+�1#�LV��Q8���jf��4����8�2������';�8��mo�kFdۼ�1U��@�c@.�'Jĵw�;-���8��z���ja�~��2���#�`i.�w|<��@�5�Ο�Ce�H}K�z#��ݛhi,mH��XA~�B{+ch���9��+���`ɿK�+��W"aE+FD�?��m�S��ӎQ6E\��ӷF��Og�
��u��@@���r�Eܬ[RM� �*[7��*#Y@h�}�Fe���8l<@���*5�����5���D/ ��|�Fٱ�w�_�i���4�F6@�En���!�@�$V]���О6pM��Άb����!�
)gC�Nȯ��1��x�� �Q{U�+~CZ 1�d|��Ze�c-b���xc�@Sf�w�Ѐ�θʘhzK*U���	�&ܘq�V��y*�؅3M��s��||r4ņx�S0d� �x�`.33O��z�NS7I핈�fȗ�B�����4"�Z�-�ZN���ʄ|��*��vֻ�2��S����A�������51�6��%�wX*{;��c�ݲ܏/�ۦ��^�[�fƤ�d�G� kĘĶq;K�Rmw�tZ�CB�ㅧ�4t�v�Z��Y��[8�L����ذ1�ʙ�2���W��L��Ϧ�7��t���S/�t��I��G5�1Z��C͹�	�<�XlxVHYEB    5f5a    1490�S��[0E�E���̩���K�BO�Q�f�n/.!J�-Өee~�W����8>+t9 ���4e��6�Fă��H�l����,���14ұ����>��&M�'��I�YJ����qվ�O�H��hed�,b�}ِ���k�o����D�1Oo����s��=�rP3�>W.D�l&]�s�v���EF��j�8�.{J�v5)��LZJ k���h�4�^"{9�O� �o�{Qa��gu*Mj�)"?��$��4��Qר�#�u @R���b��Oi ����Q#6K6I��	�#�I��t(z;�1���b��;��?$= ,��t���67�Z�h���Β�_$<v+�LR���M'���t�揸�X|Va�����ͧ���t�r��yM����n!b� ���6ɵ�ﮣ.�$ha��q뙠�D�����g��e� ��Q�Z2���G�0ݶ��f��D5��O��SJ|n.?@dUH�1����5K��h��1I!�?��â�2B�Ք�G�x���8��؛�\j�i�fXb:]�"'g���ɇ�w�')�N��+�@���5�:�� j��	Nצ�<˵�
��O㲔Ƹ�~�n�HBp�1|���t����ZOx�)�oدd2�Gl{
��I�9vHc��V?�0��X�P���/�b���2~'-q�V��h��w�6Tjta��S�*{���D�$��6
���d�Q1���ן=&ْ{��J��[�e(�dL�@��O@���R��f�ƫpA_N�t>�����IJ�C��,^����:����;��_F�k��ܼ���V��;9������7�
�E���#�%{=@�0��mP�1�����'3���#��(W����HiH�!1@��M� e|���1yِzFk�,I{[?{msڠKJsH���*@|��z�o�-:���JmD�w�۩Gmu͵��Ś��2lT��V���М��+���m�����K04�e!ry-dp���_���;s�-��zGB:O��M�t�4�u]ɾ�G\ܘ�e��,�ɨ�kv�$��EJ�(  ,�X|JS��)��m5�0��/!��8%�E0?S� �MIj*j��w�z�.��߼��p��| �?;B`;U��Ϥp�Ӈ���MF��+����eJ�0<_��jZ�M*ݚ�d��|Z�����Ξan�4�pt!U�,+�J\����f5o�vp� ��e���{�(���FM~}ܮ���g��W ��Ə�uP�kn��k�듄G�̰��#)?a`�����|ŭ��r��~�J��8�ze������ ����̒���tx�'�H���--w|�Ej�CG����<�#��ZA(�S�,�)�k��4������;i0$A�G^�M�����Tʍ{��|m6:$�����˓Ғ_>�ϵ�*8��5���7
P��y���&���Y/�QM�����N-�1!�g*]3��|��Dʋ��܎�pH��}��N� {��oRo� ��l��8��`n��������V��oLTO����<<nQ�â��d�^+����;	��yR,�]���/Mv�¬�����x������;@�R��%6jx�'�	��)���@k�9.ٝ&wϜp����g��f�ޤ5�P�+��)�փ�����?6����(����<*oCb%�8PW�C6.������rF��!ƌlϨ�s&%s�"U���
�Wh.�d�-�<S��T ��1�I�zbK����n�,������:g2-F\pW` X�t�LK�^��f�8rj�Ɂ��¢��e�|�
9d����8�����Z�;�*���D$O�����6,�,���	`~-?83@���e�z��X��1M����񇞩S�9����ԑ!�+��gk�8�B����#�B�O!�Q&^nv����g
#^�ѰǍ�]��$�M�b,��k�G�nj�݉,��,�����9�A���~�ƞ~�A�]M��~��-9M���>M?&ph[�yS�W�K��i}��Uv� ��Ȟ��d3�}@��"�o��k�c����#e%�C:�� uE�Bz�$�-�'m8��@�_W��_�.�'e�J�����*	�Á�\�#�c��l&���{���{R�=�ڼ�m2s |�l������\��X�%Z`�n�^�ǝ�)p����%���F��kv�������yB�V(��>��i��Z �?���ΑQ���}�"y_C�c�����퓊�N�I�7o�z�f|j���©�9�=��H�]C9��%�#�D(�_t]��Z"k8�B����&,������?4���ڳ�h��	��h��q8�R��W$W:\ý��R�L��h,s�ߚ�#ys묵�?טhi��}`��:Wkx�����)p&�+�M�ac�_x��傠�8���'�x�b�s�z��׾Lч2A���R�;s&)���V���yN`�sƒ�@����{�J����Y ���O���at�$M�-��3 D�m�� iy~�qr}�?l���f�������qJ� �u�CO����# �:�Q���ߖ��I��g�Q�0�-oW�w%���5a�73����x{����@t�e��$G0���$vЍ8p+z���a��P����\<�.6J}�}��[qg�R��!(����k�]#����/�y�o��a�_V�/:��AO1o��M_�:�&}��R���� pOM��nFjp��OPN�8�l6�����e��*QJ{IAp����a��Ɨ|":�8ae^���[w �$ X
���B���[���4�u�X�Bl9����m�8[#��K~���Ը�l+��q*�1���s��S)Ce���CSCbru��}O��+
.3ꎩ`�ޟL�4�Oy��CLA7�䊇�œ�b� Yr��eXc�$,E�C��$�E����!�F�����c��x3��D���a"P>�}�-��~��$B�&�VÃ���܋ۉn�G�����1T�~�9�q��Ib}	
����j}#m��
{6>�-����e�N��?����`
�f��ߗߠ�����Ihd���B�j�������\�X��}�.>�z��p�	�D��q�ت��8x�xk�&�0��%���P���9i	4KAY�5�� ��i�5�-Of���d},��2�r����ͦX�-l^"l0�"�̛@[��Ӟ����3�hd$P���0zY���8���q�e�q%Y^�����t���bnDD�59��'�6@�x�Y�U3���ۀ��O�2�V�[O�V��[�0�wq���O����u�z��x�Z�Ovk��v���wcoi�m�ۉ���ʾ�ÿ�AE�6���V�\m��l��=s�Y�]�"��"9�b������ '�߈�+�d��$�M���h�p�E�ȓ���1ZB�̦��{e�c� �9)Un�&mj�>�I ��gS�e�и���=}iz��v�p��^��1xO�s�~�~*%iӃ�b��q��(M����V���W�+��!B���4Ԑ�QedϦ�������Bpl��KtS�U��Ƴ�����<[����>��V� D`�-ev�secP9_�@�W���⇤��s/�Vt�B]Z����O��E���%"���@�s~�x߷r�n<'t�.@���q���H�.+xr���	�˯�U\�W1����0�k�-�;�o�$<ބ���v���[8����~�JK�xʗx;�0��(����F���!�h�u8J9�"�i����&��>�n3��T7E�js��3�'|��u�x+��x�Q@�8��a./�kA�NE\ěKv?l�N��;�|���9�߽����o���=]�,a�L�y����%ʘꮂ$�G��^�۸_(�a�t��u��&�ܺ[ `�(D�5�Mm�҉F�)�b�v�sU����\q�h�W���8堜*��˝]gt���v�T�?D�4!��>i�g��M�}����2�ҝB��3�^�j��%��dYL��-@<�(X�қߧ���1^�j�6�(�� S>�h�����`,��ΰ�RQ ���=��F��4���℠��np�:a�.P�PCr
�N+��T�xPo���Gj�П�YYw��Srz��<�3�HȁY4�"۝��<�$��;��!j��AI5��V�����1SP.�q[��>�� �E�� ��h�S;�;/��������H��]�� n�3��"�1�\�}{��Ť�{���[{�i�Dz�o�w�J���$����әCW�sah�A����N�L$�Z���\j��/P�§�]x�'����ۿ�#��?<@��е�7�ag�{��S���q\�4������ͳ�U�+ԓ�l:�M�{�#����УN�oHo����0�A�i[�P�`0�̛{�7(egCI?D���qI���ç6J�D�OҭJO��J�$����>+�)��>�NB3�Ih�A몹�o�J7bܸp�V�6�8��
��6��HB��EZpd.�԰�mU�}bu���p���r��`A!LY�:r6�R����U�]���[oZ���vb�.�)ow��?�r���[��;΋�J�,H|/�H��|^Ix���l��
��ˬqA�ېH��/$!�B�����DY���al���M�_f�ko�}�"������
s/u����/g�'�`��<�sN�(��X[W�d|�g���X q�^ %��n��w�q�c�A�-ʾ�;�PYH��6_�@�a6
���oɡ�qmJl�:"#ѪeJWs�T�0�-S���)��ts{\��a -ߧ�<��������e6��&��H:Z�8rJH��b݇ͩ:�{!�b�trѸ!O�k���P����� ��I��70��\	��$#�>�|v(�Ӑ����&�(;� �#H�wc����b`%#�y���2�<L��'G\�%�8R���o;����(��1�6��8=��-�5���z�lן>�	��-ݩ�rO�ӂ�hgӹGl���7�"Y�H��#:��tK�2���`��d0(��f���t� �I�!s����n���?�]'��E�xYʏ��W319ފzT��LW�{�{��u���H�E|:�@Ǆ�k��� 2�i֖��B�jw����u��X�Y�O�M/e]�M��V�\{���!�t�F�n���<K��V墀K@�)Ё��^�C�Bc��"