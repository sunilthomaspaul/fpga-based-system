XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��f�AU	[q��Ѵ�(Vi(9_ܤ�|���PÈ�("S
�SV4����3J^	#IDjyH�k�EBn�jzǸYQ@&~�x%,a��۶>-��<��o�K�� XW�wΟZ� ֳr�Q3�J�2��>Ҍ������Χ���s�j����"�m������ά=�)��i�;�ߏ�xV�"�w)`3;%��B�4��Y��R/]����p�}����1�`zK���t���s/%p6��v\"�k��
Ah�)l�."���"|X`lG���N��Dԏ�����e��x��/�[��&I�[��CJa�ui����Z(N4L����o���fx),E��g���,�A��@��n̎�@>2��.R4Ԕ�}���5�?EC���`�o�'�����#q;�F�˱�I�*���Q��岥�4�<�����^9FZZ>��A=&<��~Nn�M�>A�����d�,���@��b,h�C�uu'�CT�C�����F�<Xe��t93���΁����w0Trڱiq��O�|�	#��L�m�9`��J���vz�E�A��dc��M/�uIWN�0�n���1�ӎy#���׮ɨ�6;:���)����K���\���]`%D�o����{�"���n�^]xI��չ4�R�7�P�D�ŷL��ݮ��Ӽ�'n�/?�VM�3�k~��K��U2��uF��
Y|�H���HT/?�b
T�(�����2(]<@�E�T��J� �Ѣ2�oυ��XlxVHYEB    159e     7e0<�C�<>�0q}k�{QS]�r^����Z	SL�&���퇼��\�*Ft,�mܜo�~�խ֫V�_:��L؅���]q�0�'f�<7?ǅI���&<^��9���Տ��5X��ᖋ(��rY���9���\&���^��KC�������Rz{� �a��߅�a�x[ܧ�r�9p�a�#�v��ds�7W�Q�G��t�c4L���Ql9X[x��A�i�
S��ѧ�+ʮ���y�hZ&�cG��>�VS"�䳼|5Ob�O. 3�
{�4���O:"<��wwt3��M���T�r�a�9��U �88��j=�۸���|(}�� �ر����ܨs�t�%)�<����i_I�Z��a�'J.�w��71���& E�2�.I���d�N�k��O���i�5\���,c�Q���S�rx^h��x-�=J+�`.�e:A�us,��ݍ�@cc��%�l�38l!�-`l,g�7���R9�m*��
�Mp�RO�WS;W�zy��,x�e!o_���c��`������C��?�Dc�ճ��,&���!O�+��29S�LU�����G�%�aҘ�¤�S�8Ui`᳢��p'��\A��kgd��
^k��4ҕǔ�8�X�����	�뗐x��Z�~�&-���d�f��n��a`�������n�;9ëض�k��l?{�{g��P|���W�/�/�P0�8��	ɸ �^�y�b*�߉{>�$k{��`]���=k&W3��&$u�Æzt�����q�3jN���ԥ#p=XD��\g��D�?��Ĥ��11A���F�mIWO	�d>�L������+mV��W���&�J��}(���:��w�b#��#N�`�{
5�j*;�e;��x����Sw�v�k����)�ϧ��'m��v�9>�\�&l[�h�T$��"��mϬZ�������7������e ���rlU�/.atV���N�k=8�=0�^��)��Ȱ�K2z����m�*V��AjL7�w�oI�Y�Bs,���o������X��[�q+��'��R[�O�'|��\�"���d�֭��E'��`9��Ԯ�@�"?0���c�;�_��kt(�!��*[����w!-��J��LNs�f ��#PA3-?m�XP��m�Unx�K��}�K��%��K]s�������,��v�?Crk����|7&���nb���K�?g�UF��[�J�Z.�v��F���ٮ�Gҥ����UO,Ċ�c6ኾ���Lg���hZl!E�<⹄v���K�7�\\C�k��w�*�Wj`MN��6s�B#iF!m;d(-~7�J�7N3i9� �.��YP�:�
z<F�:�6��l�M�쨺 =Z�����ם�n����l'c��F�d�������@��G��J���d�@(z:�,6Z��%�j{�+�8�f�f,�y�C��=%�������_s��	*X�<��kϲL��~=��WJ���b�.��.�͡�0(`�pן�FBG��yr�#%<]KփV<�
�c��1ʄ�4r��5Mx+>��GIg'V
�+�_By��8^����6�[�m.�=uH! ����Fc>��i�$����/vHC'�X��?1�M�?�^b���9Wu��LW)��A�yH�ߐ�����;qz�l&36�|�a��!�߳��Βd)w�-�/�7s�c�Ҹ�$�;)π:;N<-v���҈}�@�/q�� �{��Z �j�~ֻڿ!.���f�x�������:�>}Е�L*K����$vPr*a��X��T������(J���Cnζ��P�k�����z�H��f��Hw�ݐx��h��-��&�
 ��+��Xz���z�HЗ�.�$[����*6�|�|�O)��P�!��m�e �DmcK=1���.����.25�>XH�=�T�}��Y�O�妿� �!u�)�zL���V�
�p=/%TG�����'2w��+S8Syf�j
fx����