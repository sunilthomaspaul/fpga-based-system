XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��gh=\�Y���Cґ����r�zI��m]K=$��ӵ:)I
a��e�`D(~Vm�6�1Pkԡ�m@M]7	h-W�� ��(z8&������6(�CC*����~��`�?� .�4Ɗmҥ�\���w���>.��K���[UUP-�_tƞ��"�6ʶ/Jx81�ҳ��Σt��y�H���_{����X* j~\-8q��6�߈T�Yd�b?ie�*�����y�=/��8?�f�5`�w-p�������u~��.g�G���t]��ҎL�;w���Z��J�� jވ��Ƭ#���؏��rP.3�G��R5e�����2���C�}(<D]x�2O@Y(�������C^�5��Ώ_�2ڏ��G�Q_������M#�h��N�mC�b%��Y\���o�w�
g�^�L���$�a8���Fcn?�0U����4&���n�V�$��D#
�=l�&[� �~���0�J�����g�x+�(e�����������l�;	p��f�c2�s�l�"^`�n
�u�`�
h�=f^�\jD���\��v>'��Q��}y @1�#.��@��dG5�fgJfU6�W�9Z,̞^�l�Rk�@�tC���4�e�!���\��iWx8��{R�=���E�'%#������mS�
��6�<����&�3���;7D��l��u�)���)�����W�K�E���L��rhK`�tj@S�O�
�{Ԟ�|��uoz��p]_���i��XlxVHYEB    118c     6d0���zc�.�&��䨸��x%X0��\.�����+�(����R���b_~������a�7Rө���o!uP"Mw�'�60�������?'y���d9&���%cr�����v�MG�.������-&I�ݽ��t�Y���*,P�AO9��QGr�p�mCNWjt��Y���6���5T�w�}8����'1�'��ɿ �]��G��5)FH�~ F���F��}ⳮB0�!mx�.�E�\+�eBj�?ŰVċZ8bd�%�"(ŢB���JS82���+2���w�W�!����/v��m?��W�gݿ=��l�v=�cn}@��M_E�y�`sK��^Nb�Q=�a��v;�h��#��5Y<��NGazgoi"F�x��[_���)[ �	�xz���\n���Re�D�X��g�HVIF#�P*z�����^o3+U�\#�ДC�=2u���r�D��mm��\A8Ԑ�u��&ݜ#yg��@���M}=ֹ�Pm�lˮE�Y/���h��E��+��ͯ)��l���֧pMs��K+�����57s�J���"���<���TAkj�%hp� �Ӥ���Q�ߛ�쇀��b]��3IMB�h��s��s�����
�� ��GΖ��_�*��1�%��o`!v`	����j1�26��9���'��p�km��}2��s���� 
#U��\��������L�+\Ǯ�f���Ykb��ZR"�>A{���7W�)Jɉ2���ZrB2X5E��=�BK|y99\x����̆5Q��Y�.�lۛ�ni�g�*	�`�A�RזO�  �I�G�f�qGk�֟o�,~
0�K��6����ԫ�:&蒩���h���o�S=�����7[�~�@z��V������C�ǎQ��3�uFwW�7$�7�q����:n��4k�e[Ez9�@��� 4Z������Q��)��͎V���Li�Ӌ-G���6;8KZ(j*���\���Ǻh�����<E��ϮEE
@���~7x�H֓t`��e^���/*�_��>��f���$Kd�d��U����ػ����$�B=P����ٔB�*?i��Cux�i�ݐǓ�?��w�N�"�l&ކ�l�A(ڟ+���د�6TIˋ�2!D;r��y��<j�ۜ�����x��*eʘ�r�J��{�8�Q#��C� n���]^��>��C�S,pP��#L�k,t1���J��Ir'�rM,��+��zI^:�&�"O��E���%m�x��a�T[��+Sj$qK!�c����.GI��@��'������'4%��lG.��u���W���q��	����E��a��luh bXf��tZ{���"�	oN������9ٝ�97Ղ��W�6�F�@~4�m]��`,V��%�/�$0��z�̀XԮ�(�I7X��]�P�z��:�㥚���~yb�Il>�b�NY�ZM�-_ߪ,K�T�6�r2_q	�_siBD���㽔H|s܇	��$#��-ю��?�"y�T��P���%�	i&|��N�~P�r�a:��)Fl��.�v�ɰ���&cK)&϶�u<[(d�JI�I�Q]Y�,�"���4�����n]$��=С2�s3ê����p�H0z *t걠LjC0�~��u
����5UXQ��h!��.8��&�J2�(�FH.+��pƸ&+�ނC؍­Y�Y�j= Ba?�L#Т�߸Ԑ�q0