XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���ǉ�z��N2��#�YGb:�W����`&���o@3=�����)J�}�*�q����lvʴ�~�_�A��[@�"牄֑J2�N�~�ɕz��G��ɓ[;�b�3�`YB�y?�	�4�>����]k��)���f�㓋$�, PA����N_G!����������.a�Sq�-�t{�� o�uޱZ��X�{�Q���`��y�kֱ� d�;.ER��NFL�l�ښ��BDaw��,[��Ϟ�v��[�H����6������z���D�w�h����H�#��Fc�f�*�0]�|�-��!�עe=���N�(`y�K��p�o�¥�?z����]:kr�� 5^���ҋ�qn3ǀ	$'��QK�ﱚ,J��RVnޛ>;�;�� �Y���:��F��Y顏59$�|�P��E����4�^4����8��i�-��y[��no����n8ul���������6GR���Q-��k(t����w�u��v��w
�K�!\�Q6]�H�/�1���N��z��}_��$�R�غ�w�+�E���X(����ש�'}Xv��W��] �Y��q/]@����M �xW� �
Z!�=�l<�.��B�A7��1�(eO�l]��v�֕���I���w(T�)U͖�c�Z���+��e��ѿ�	;��'v�K;!n��G�Td)�˒^ϊ	�E���[W�h�̙�p﷾�o�����S6�{P
�ѣ*�\��3��S]�n8���:XlxVHYEB    9653    1860�KX��-;��\g����E?��-\���^Q.gUTB��7�]�(r��臝^�wH���usu������(Q%���&�x@��y0cND�}��ǒ�x�pYރ\U*A�� �A��]"'DE����ϋ�L5��l�{�~?T�}�8[�`�����5�43�!a��~7�l��^G8C���ٿŀ��z��<򆮣��Ν�1��ؔG�)�g^�$F�m�
�Ra�	�ε�!D.���af�L6�4�؍�ßmy_-��a�\�MX5bf�{k�pk/-��KZ��փ+��C�5vѬ�d�_6e��=@��>�������+H�%=�������cjp*��E����|�F��axw<��ү�}�M��~� �O�����~�5ҩ�b�`��{?S�F���+�~� ��-��!�i��r��P� �>`�-1^��Ì���>�B��_�ǃzŶ������`�m����vBB���[P2ث�a"/K:fZ�0���\���$	>�KS="8�+]qQ\Z�Q��Q����c�!�ަΎt�T�Ҙ+�@��}b5-��H4L��������ih+scv���}�E�4�XI6�m�P��p7 p�����Fc�w� ˳O�
^#������"�X4�V���+�q��6n��˾�h�R'|.׵F��t���X�z	n���¼�$d��=UW�M'���L��f��D�"c�h�.`��9~:¿ե\��*JGm�������۩�d��:���8|��qa�/L��ID2�cTݹY5
~�*
�^޹ �/��+��t@��d��Q1�i�$����eW�h8��^��XG��ff��RV&;W}��^x��x�"��I�V���^)�ά�<R$�xt��5O_�[IPCV
���ze���JRh�|�6# k1�7aX���@�𸽬x�@�>�jكJMA}*��\����??���ɖ8� ����r�`C�0#��^�MBg(�b����_����%@�����I`��!W{��K�W����8y�S�>'�8Ŏw�7��M�)�±�Zhꈴ"�]��[����X���[ے����$<���([|ݻ�	�>hhմg-�q�`]�q^��:�ϵ���`&��\]:��"9� ����=�:��9�6�d ��_�g���s����<�J�g����л֧�����B>,�K����-��D�hƴ��w�dV�ب�!�X{Q`���1��So�,�	�G0���a�(I�~y�Z����E+��-�f���	�Ї�Q�B�3������
�yĨY۬�8��}�5�����}~�)Fg㷀9^�0e8����TM`�v��M���	�sˀ��qt	�7�j'^; i�e���S�@��B�,\����&��,B�@�A�TD��b>'�_2%�8Y����2���L��x8�k*a���g{a��Ez�J�t7��� ����i�3�� Xw���[#&}��������(�m2�+w����u�%�K���P�H%31S<�����Ԓ0v;�̢�ay�����x��_:[b
Q�����e��7+��sN�)��`|�Qg����<i�"��������~#����]�.P+D���Ѹ��pN7k��g�d6�͢��.�U�1�����p�*.�v;�'蓽epB4�� �Իf��Q"	��5'��~4��񓾑kZ��ܸ=�]ӑ��YC��j�Ov�5��ʬ��7*$a��m܋� ���2�KeEC@��z��Ӫ.�Մ���$U�m�}ܩ��_sl<��A���La�_xoGb;�'�Q������6Y+��5��	�ϙ��n|�,�[y�z���J�I��Zq����;IZ;���!�a��+�Q�:, �����L���"=%�ٵ������w�c��_aѽ�T���_|r2�)x�E����a	�`}d��$+Ω�h�f�P��`���ٷ,F=~>J�Б| 8���[� T�z�
Eb0�9��Θ�v� �V"q�f>�R��=j.�Rn3��t�(}���S�^	�8�1��F�!}�2�5<Hn��y�
��]~U.(�e����O�SV��p�*��Z����X�a��Lҽ�������X��5�J��bK%(�^ٻI��b.�z��f3�m���24���M0yCFc�50+b���ٌT�(� ��f:۾|b��`l�
d��\�;�#	6<p�C)��YN����Έ焩���P�{JD��H��Tg�f�b�#S�-��+켩mt����4����Y,�bi;M�ZM�4�j��̦eVMN�d�8��w[H�������~�3�&XCk���Sgk>4�՗�tE*�\�O�c����F7�ؙ+��d��9��(���H��N�ߙ�.H�����<4�+Ȃ(�{j�F|[M �"��9P�����Π�=�x��Rg�`�����5��Ji��9��0D��P�^��:�!�!PzGs��T�	b������Dt����p���g��Y��^ֱq�l%��b�A��K�.��n��Х
�ȩB���
�
��gzd�������<�=&Y�7v�qzF�[G�5�,QPY7��f9m�I֞�TŦV�յ=mL.T��$���g���y&%�w�p`�n��8	�(ٽڷt�r�jG!٤}e�Z�D>7�p�2\� *D�С�l@⃺qB�_Jr/#�U�\X���1S��T�g\I�٤e?��.��U��J}ªn�T�9G��ۙ��^�����)<SL��n�#F����.tH����"��Xɦ�8�Mi����u�n]���$X�S�?���##�a��G�c#V�pUl�qr��$��o��a߃i���֌I������p��W�� w:��j�|(NX{�_��ޭ6��?h`�cG�nr���k���7�����7XzYǉ6q�K��Nmd�	�Ǝ��v�����-�<s,Z��L�R��';���u�5F�r��R�cS*sOo��?Q���츟��O�l����Ɗ#��]�@Ft�%hڄx��Q�'�ЂJY;���D�Q�jB��\Ǜ,�7W\��˭�-UY�]j��1�x�R>?��=dI��#��svy�߮�BD��Sq����t�dee���c۴�������%�\��p�F��i\vb!|ʥ�D��|�Ө9����γ�~��ٽ(�0!U�&�F�V��*�@��4׹�"Պ�!X9�f��:��X��A~g/ҁ�W����gԥ*��b%�B�dG|���aV�z�nq�V�C"k�����T%qx�`��D�g�O���GYj��Ų����hd�;���2��_�2x#x�9n��q�bU9����?�;/"�Z�����?�^J�f7���0 �2S���7b��_7��4�f���}�ȯN6��B�������'����OV�ibr�Й�7c�!�XX��*�,�Qi�3��?����>�����>q����o�툐�(��{�+�{([މ����/�/��W���ǋU�?�k�������_(I�4�����5�'���ڗ2<s�It�'���>�I�ĥPO_�N�C�^Cꟁ[HAa��_2��L�`L��;ڝ�æ�byS���w��D�<�.'�%�P)�Ç��������P����b�p\�hH�rn.* ��?a��5W�{W6t�w��죜|���m���dʐݐ��@u�-�U�&LI{̈��'kq_�Gx�o����P1���AYX����*9�����c�̒w���|3�$-���ZM+�>�b�1�Ӧ)����\f۽�X����ߣ�Ƶ���{wu��i�ɭ�+M_n"���"]K52��N�W����G�	]��}2u�]ݒ��A8��G�{�7�l��S�2=�?#dD��nU,u��n�dK���n��m0���*�Z�>Y�߽��ʵfyU{�����������,���X��&V��5�*�S!��UL�{	�����Y/�f�'�c%��`�q(��.�c��]tp��-�K�����0�j���I������"J9i|(Jw��u�F��ZVX��=$���b,P�A�\�½�����C��4I� ^V�!VUL\���aG�� 2��� ��n��7��xI0�IGb��虞
Gg���a曹?Z2�1��{�W��"�!�=�P��q�"eCԫ�&��"a�D�9q���˂�ژ9��[��H�f���_�N`zK9\���bfډ_�s��f.��+!�l�#1I&w(����ƫ� !2£t.<U���@��"����I�����/D�!�x���a8�4�8�89�W��HC�	#ATB���1�3 q
,}IO��=ՠ��&P�a�\�@ׅ�������n�ƇbB�<����5�6pc�tC������,��^����~o6��ja�2�'��¦)�YcH�\�h����\���m{�BŪ_���㓣C�u�~*�1qi�����#A:��<x��Z���W8:� ����ʳ���F��^:W �

�<م� $^	�	�Z��9�HG�#)�^(�4�N$�͘�_c{��oc����A���Ո	tx���LZjS>9�,`�6����cn^���5=:��R)l��[����>�k�h�=����E�����oo�('T��ƾ��Lh�x')���m�@̃��	w�O���U)�qLy����Kp�{��	^/1J<�q�*j�gA6�I �`Q����gw�?]����q�M+ȴ�3�3�Ah$;˲է��	&��k������';�� ^^>=Z������7�y��i[	D�����))k�!��_�T ��GF1Ñ.<��j����D��W
�S]	�����?P��G0�ë}!kS�,�uv���M�v��c��@q�tѺ[c�0��$	Me"����*���tk���W��#�s�q�L��eKI�H�\ s�Q��0��u���~@���r��˂��k�FE!ߥ~{�+
(����7��'-u�+�/�-z&�H��͈���?�4���(���ˮ��A�|�Դ;w��mSg��r��>y���ɻ�ޕ��c`L�E�ג(��dlE��c�H��������o���Yz��ݟ!��P���ɴD� �I��¢B�G� �͉������a}$�a����H�r���%fqU��yd�%��"ü�I?sNs�a{O������06�I���eH>�4��%�9������c��\�7�i�ȱd$^{n���u)7��yܟ���Ok�좨*��OJ`�wQ��ÔBr�ͼ��r��8Nhh���:�.�¾�)��I�ڝ�@9�ó�|V@�AH��U��/�J#�@�$_�x�=\��P����x��������ñ�p�b��'��(K
��36؝�M�-����C��[�����D�]wT���e��`�R-��*�T�z:>�F��c���6��<X���JR9� Jq�5������_�$Nĵ��au{Z��O������h�[����xt�J!��/jTih��X��7$����u�p����i�&��}�w8��Q�\V�چ1�h.cy�N�Ѹ��Y��`aP����B�9�Za����=��m	�{�ʋu��#6�t_�����B��B�ȎT��~��<�D����_I	�Kۃ��h(��Q!���,���`4��Skxϟ�Q�ɥ b'UD�d�D05�Tpu��$��25Qu*�"X>p
������m�
�	C/�p��4�=��ߥxsn�V�N�1�N��h������$�	� 7��h���[����WoA�3�Ps�`%gI�#>4o3�v�>�}k�9vl�䎪��9Ϟ�i�eZ�r�tJ~T0H�C*D�  ��]}�_�KoH�N&&�����D�ze��
��ݾ���M��m8<�%sW1��<�Z=�Bs��������36���Rڧrd��P�Z��6mP�Л�Lݬ�lV}�U-��So�"���8J@<PAh�����I�>t��zIǜSJڝ٣{�j��u�|yG��b�j-�$��V��y��H9�0m\�)��#}K`�ګ�:&�w���v�{p�"�h$R�gl�G9ScȚx.�d�>�:ΰ����>.��uGf�����J�C��8�7�M�����w�c�I@N�P]Y��ǺM�e�$o���,���m���