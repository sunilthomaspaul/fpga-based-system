XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��º�y�Y��'coZ��C" ��w�B{�^;�T��!L)�
훼�����a�*���?7�f��M]����:B����Ae�m�Pyy�U�4�F#f�#Tݚ05��f4]�(T��n�' $���+��'�8��R�lq� �ˤ�اO�	����?��-�$�[�5\��9>�Z����"��{dɽ3��t�Pe����I2ϹCU�])���� o�0N�8��NP	B �:����=�`�Qv�ۡe�7?�������߾ѥ�*(�$���>L���BoG.�[�7]�$�h"f���͉!�Pw����/��w���Uˠ/�P
��#����.,�0\!&�&�#���n�Y�M�B�+O�xQ��gˌ�o�����x�����M�����74�CP���T+�����M����0����m^�T�J�'f��g㌟�=Cl��6'���=+(��X �/��#�m�q>�6s8B"]��P'��d�+��Ņn�"�k����	���G�Cl�T�����	$�����bq~��#L�'V�� *4��8ױ\Gʉc��⾈����k)Ss����c�]a�k��V���B#k:�m�l���%�?K�I����T^#bZC���F�$��)���s�X��Y��}��r�NS��ň�������Da�P��9���}�ۦ�ϣ��k�1��/�}Pr�ki>^d����̇B��
R>O���n��H�ջ�ŀL�$!�L�j�%���!�kxɛ6�V�FI(k�XlxVHYEB    4071     db0軞'%���s�y��MP؎_����\SUV.ⱈ���#��.A�^��I����2�:{��]�o^�g��mn�X7+�>�[2{�ۧ��-U��=IA�ST�B������]��Y%c���׳��ؒ�vO��[VH���
�Č�$��Mx�	��<'D���u��W��a�w�~'�J��|x��H���ϫ:{�Pt��M��B_�+rp�Ԃ���xF�����tN��/� ���Pf%�Z�v8��ά�8P���Ϗ��\����K���C9�ŀ��h(}�|�E*�\4S]F)�Ij�IH�����*R�v_�k��r4!7ʏ����]W�tU~�Ү�헲$A�����4�n�5/�5-���N"�=ufcv�]��D)XS[xԫC���Fw�q햱ܫw#E?ݎ�/����&����ޢp���T���8�;L fۣEȫ!�t�R~�,]��CYvV��d����'xs���SA��f�W��#�
�T'�&�|DoNC�W�>	
���9�s���ࠪ�{wMI�ʋ"@�%�����~���Z�}�~R���R �ϊ�JA��i!tB�5��0q�椌�<����y�gR�Smd>=nTr�"��i�.��|o�7��i�����P��P���v!���-Q�^��{Ar2��IɈ6(��9梏G���Q�kb"�����SG_�p��ܱB�sO��'��s\��L?)��.�B��Q�3��v���91O�KB�#*�ֻ%�דYO�P5`��L�@?�(콨z�K��ݣw�V���J�$,x4Q�R�K�Ih�Q�ƣ���"D�D�ۂ���;�9�K4S:��(H�w�Ƨ�A�hʲۉ|cN�z)DU���E �[�.�I�鲅T�zi�l�C��9r�����\#��KdK�W;K|�g%o [�I���{���Y��R��u-Y���*Ua�o�z�o�"6}�Co��yχ�̈�1,f#'�r(�p4�"�0	�8Ft��zT`x��hf��ʌO	��e�8߃}�#¾οu�|\�� ��J�H`$Hr:ۈ�LT�??���w�c��͐�X��~��|������W�"�c���HK��������Y[`J�-�54[�E+ݢ��#V���nc�t�V?����V
Q�;�{P�����єl��7��ˀsﾆд�A�j\�`�`�-+{G?\�8~���H;�Ԥ*��{��սw�mg����m)�f_�CΑBw�Gu�
u�r��Ԋ�!���$K'Ͽ�:�rKQă9���nV\9uN��\���W����:��+�*��#2T��U�Y��������Q6ގ��Ú��
>I�Y����?4�ݩ*���d����-�yDb��͙݅�8�������Zf�od���g#�!���2��>m����/��".�s�\[ 1�9���bR�ضKl �IN(#���G_��0I���ڏ]���8�����moBq@��JM_�Hگ*�]Y������%�`[���H�z��8�v'RA�#`yq�<u�~V����Wgz�{e�mӉ;]�n�֋T̖�ȼ>*�+#nI����>�eb��kCd?�;|s1M�9ڹK��Vx��J��h:>�����|<��V�?u/���5�#�m3q������H=� �gz"I4Č����l�8aM!�Ս�Y%3j1�=�̥#G��+O�l�yB�i�(�I�fȏ6�0f lj�.$!�fS��K]+�";���Е~d�D���O�՜	ua��1�U��6�u��������K��R�΅W|��Ͻ���-�E?A� ����z�������"R�x�]LCzyO2Ƿ��w�	�r�sn��M��>�'��c�v.����O�L�,�(y�gRa1눧�Zi�[K	����6=��:S��h�o�ϕwZ%��9�������Ȟ�R�荕���F�X�hX�Iݿ��mC���~��8)v����	>��0x���A�ifIm��� �W�)���/�1�3��+�7�����6Ӗ��U�� �bM�.@z�.*�:b�K}����aȊ�s����z���4G��F�S0T�Y���O:����H�D�_�o:d��_A\n��&\|w3|� �hPi�\��Ӧ�a]��bچ���Q�;�J�ݖ)��ҥ��>g6s=Z���$?��#�x4�2�v�Q��XǮ����iNqujv��ٶ�r0���7a[5]��*Z*)AV����9H&��8p!Ȯ!���(]�D�Òêc';�A� G:R?e�4�j�#��aڏ�B,{���E;6*��l��P?	�F~�z�k~��r��Jh��&_��I�Yj�}u�G١zz�n&k���X�͖�P��]�U���#,H�n�(@���؋�+R���S��t��rAL~
����2�ml�|�z�WH3��t�)Uj�*7�Ce)H�\�MB�w�v��D��9��@�RaL�D>�|`0�载H�����>|��^T�}(�6����˻�'T�de)�JkM��>�?:?I�(�f��m�]dHJ7/�c�@�˰�K]����خ��Îj����>��ZjϢ����Hۑ�����9Z��kFW��ncT,ಿ���DEʩT��-Z'�5�����0�z�;kg��)c�|��|W�g��"zQ�M�%jT��{8,$Gqѐ
s1�ۈ��i����>��'*��a�i���"�6u*Vq,W�o�4�PXS�s�j��^,��϶�'�B���� f���@�͚P���ї��"�Ć������!�lTe�� !of���E�a�旡#pJ�A$����-4d��놃����;c�$3ZF��G%c'��K�HK�3��p%G�鶴3�?��p����F+�����{�(�0������z��`��I�P&�)�0ԋ������f�Ճ�g��lw`ׅD�kEK�m��Me\��j��YlW�˧%�z b�1�P.tj~�_4��k��̫<]��
z��M���R��p��B%���5�+9cr����Rh��-Ot-����snE�TT5��	�֕I~�Ak�j�� ��[R��\Ӥ�3����v�կ��k ���d���I�o����g<Z*yp�C(���E�>[�o���	�pws&� �Z$��G��;��>�R�� ��f�;Gf�Nĳ�u$&���,\������HρC�D���J'�������H���E�L�l�u����-5���j��w����׊rpv�����:S��e��(�4��DT�bp-�Ǉ|ƚ��C_GD" ��;��Cj hN&��i�
���	�py�4���7|Z��$g<?�N
�|/�țp���̓|��}�뿃U~T+I���#SD<���k��?ȨeŪa���Cr�3��\.�x��� )`�iK��e�)q��8I�z��M`{�S�Ne̺"��y^B'9$
A=