XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���]�*<m�o�ۣ
l�R}���S�얹�F�=�JV�SY���O_�򮐐�=��ל{E�|�j�����$^n+A�]y:sV��8k�D*^�Ƣ׻f�ǡwG���q��I��W�!�6'�����'mc{8֣��#�U����;��-!?��Á����U�������Op�����R
��G^���㵱�@Ao������p��[B����l�+G�߅���lߖ������>�h��B�;^��4�xl��~��e|�j��`=�'�Q��osN��������v��փ�f��-�f�f!
��u����c�ᲝL'o��a�>��Ȁ�ˮ�{Vs�نE��,an�5���"�f�P��P���?B��'���<���h!����)��w"�1�V�&sͥ �"�Г�6�X��pr��#?z�_iP���9�#n�?��ᡩ����O�V�&�pD��Z)t�FS0`�D��R�MR��Cz��W�_��iK��:s5KKK[~łu)^��������(&���I�G�������[�+�AU�{F�0���2��׋�6׾.�o�0�����>�7��T�C"��5Ы�/C�U�t�ۉW��o=3-h1�U)��Y1��\ď�7�k�4j��*c�dj�8���[z����;x&&з�QP��}@�"�_���e�y|9
jx/sYC8�_Y;W󬧭����'���ȴ[��IȨw��]��q�U�غ�H����ѫ����Y@�=����Z,�XlxVHYEB    3e0e    1150�1B��("�	��( ���@����e���l:�k}h�up�P,�s!qû&,~��Hp����v�k#(jD��9]�0H���p�f��C
-�tY`���?[n�u�α}u�X=�ԯ�H�s)m
�"��u��R��{���|q4�=`R�s������.V�?/a �?@���/��ͥ��8�����-�d�޹-�#�w��(�uԟ�i�Y�>�^Ymq��9xhޱMAq�?ኦg}nu� �0�S�o'M�}ʌP3�\�j������V�+�y��S={�����UQdo���+f�4�ο�"�� w+|!qN�� IH��0�^v�ÊG�ջ ��X�+���0�?�񾀉9�ɩ` Jz6��Npa����� �5��.\ ���MF��g;θ&go���ۓ�e��.���k�E�Sk�ȟh����m����۶��*)(
��R�[[�6jL{/������z2�0Y,W�ڝ��^�aGY(	o(����Ê(qj�>��7�t-�CN��䍙����0V��(}���A�r�gei�\&�/c�w�0X���P�m��;����5L�I\��p��@@`|ð�2���
�
��$㑚��4���e�68;\�v�-�8|0
z�Ƣ����Ζ��J�'�-�f�ZJ��M��� $4����Ks�,&����.���������Џ��Ycf��q�G0��pf����{�U��#�dʬNb�;^:��#G�2 ��5H)0�׮��9�t���E^2�OH�*A��:^�"z��~"}c��qL/�ӈ�5B"�q�� }Z�:y��`���گ���b�TQ�~�4���$��m�s۠!�	-d� ��T=2��%�d��'�S��ˈ��څ����p2��@���繱-j�&{Q��mf�Su��YI��#U2f_�	�%�-��������x��`�2���h�I�/��I������S�䨥���8��	�3݄�A_"Uc��HC���g���<Z��%+����Cy����Q[cBc�b�U႘k�n�ϝe��Қ���+?2̈́S��]���������Ϣ��t���S�G�iO~}�W~g�t�|�A�),R�`d��%`��01a����L%X�Щ#面����x����9�qG>��� E�-ɇ���u=w�.bM"��ٟ� �VK�f�^�6T3�(�/��
�*J�y�?G����)`�BeՓ��
�8��=Y*FI�~��T-�����C߼O}�b�b�h$�����W��4'h&�̋-��XbkS�P�@�nB�Ym���o����Zf�(zQAS�Yq�GP{���N��Ϫ�"Rߏ�ff3���'�QI%�i�����
h��-x�%S�ʽ> ��MA�?Eڧ18�Uu�� /�����/y����^�	�}X�Z��V�^B5v^
k���t�]�ʹB�_w��c�aq�7t�Tb�'N�R����2v<~1���C@�6T��@�q��<���A��.V�)�n��A�0��=�V>进K���
x��(�2N��lD�i#�Ŕݩ�8�\���f�C�kYJ��U�~"5맳�N�н�F���OkηH�2�U�T^fv��������	5�3�#�m��h�J|������k�߱�p��:�9�B;�l5:�ǜٸ׏+p���}Vאe�.ne��l�2�(g�8�70l���\ y����\x��h�^�<z.�2���dV�vu�� �&z��S�O�����w2X��3ES�v�֌����.�1]���u�'�_'Y���>}u�s����cc�!����h���RHAQ��=����I��j��\j�����o_׍e!D@/؊���*XG�{�*D>��l\N{�+;c�_	o��Ufz�ެR��<�������Pc�Q����#��, ����Ҙ�6��pX�y;kǨP83��,���B���Gr2�k�
!k|�S�<���{�
$2(1M�	�僖{$�y���@��o}UF��!�P���{��Vq���y����OX��K�p�A@:��H��n�	@���F�Cz<�#�ʴ����}V��$ޭ�Y��0��F&_6$*[1�P(3WI�IQ���ٞ�o�W���m'v�/dM��Pg��b0�e+�F�Q���-UHnE�y����O�=�DM5�� ��4�/���i�Ⲉ����9�*B:�[�[�2� �����#P�Z��T���?��ڰ#���w�z8d<�Ӟ�
�`YFH��*����5���fO<��@.�eƍ��$����$j6�Mi]~]�t��ҩ���*�{�l:�!F�hW�K6i�ť���}����v��
�\'�\!���ҧ
��x� {���ߞ��Zu 9l����
�#�(����7��0e|�P�.݈�P<S��l�H������^frI�J�^���_����1�K$uc�6?m4KXdt��嶘�_�f D/RA�f�~�mO��À����2�}�@�ސ�\WM�+S������_�F����$^����� �#,����t�1�c:�� ��̴W���4�x����>��r���Z��³�P3���Ϧ��ɘ�nWL�ļ�0��~���X�oa��F�$�4�_:ޣiA�_��2�m����	��P'�uy1(χ����H�?_Mp;QR%�5"^5���8�Abw�1#��</�؋��׿�)��R�I��uݟ�o +��e����>��K]d������?����_ˌP�^!�Ǔ���2���pc��΄�ƈ�r ��%q3�lʲh]�]e�d+���ձ�D'0�1/]Jǧڽ�4��=n���ś"e8=L��m��ĝ�l�kU�RВa�@9����w�3jf�>�n�s���ۑJp$��ܞ�/U�@@o:��N,7����l{)q��3cx2�W�aL{B�}�6��U�I��ǫ�� x[�PӲ[B<?!�:NS>['� ��v[J|9_��k<�H?Ï�?�0{�n�S�7o*�����)�J)*�gvԖc�	1��� B��־V"��i�cup{4��x�/���Fi(ڨ/n�ȷ��$� ;Buڗ��F��"h���#;%����v�q1�X��'���a
t��>�U.��&�#�
��nf�6����f�2�S#�X[���C=PX�V,4���A���ʵ��s!σ���7?�����SƗ<E�jl�:g�Z��J�a0F?	��:˖���)� ��hy5�B�n
�ȌÎ��T�:����������!Rr��]�GbtH`*�eq)�7G?x%���4e�!D}�`2�~ό@PDy�����rW[叻]�L�nU�X�|�u��b�
(��-����I��ꁂ��Ğ>��]~���(�k)y�,6�(X�6'0Ґ{�hT��������2���d\��-q����a*
Wj���P,�Y��m�:�34��f@M�h��RQ|����:t�����W�i�)?�I)Q9"/��U�cl������~�P�Z�nm|P?�݁�'P��������<����{�`n����tŤ;JrX2^\#�w 'f!�݂.��-۳XSͷ_w	��s甑d����L����l܀,l�Q�\Ƽ;�{���v`��8����: �,�K0/�c�9��ɳ�C�a�` �>-�����WN�h.�b
=�\���i�m=�~_�x��ǾP17oѝhIzA�
HH�$r\=t>�yong2M��P��$��O��*��ۮ�8�,=Ϲެ ��K�^��6#�w�6��۸Y���?Ki��%߲���8�t}/e=�$R3��&rF�d��̣QX2\o��A����P�bj�U�+z��7�!�]���-2;M��������،�Ut�!`|�5V0_1�̠Y6��R�k܇��^��#���M��'!�O��dϟZ���U��@��[׹���`���>��=���&�̫�_�vL��ouUq��2¢';�#Y*�m��Ce���4}�7����"4!�!�t��&SD_Җ3=n�U���2�2���If��=�ؓ�l�C�~FZ*�#v{�9GJ�T��ó�I��ƭ�{b����y����N���o2f�)Gۥ����,�3ߜl����Iae ��),.�@�O�W�G�Om�X���w�UJ�G=��7nаL����o��t玷�k��o	*��V��K��Tp�d+s�~�`�L�_]Ӽ$�7�Șҝ��ay��l�b�(���A��9LH�ӄD�Aygg�'��a|:���?�(Ӵ~Xo�So�p����tR���l�Q�J�:_%n`�k��y�,���ܛ��ٯ���E�Tދ��g9ʹv�Y�v�	׉.�0t<hG�9'�P�hIz�ځ�e�g���+Y���v�ܝe�B[K0�e