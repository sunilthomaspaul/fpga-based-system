XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���F�c��Z�_��L�JJ�©�-d�/��3Jk3L�P&�9�^	���R�`gm-F��V~�Qx���dz&����l�j�4ۡga����c{����џ�����O�1�J�^���.��G��m�`q\�o(�Z\��l�#!ؙa���s;���{��ϗ�	��غ��ٵ����z����؃����|NT0�P�=	�Ǵ��&�#����Ja0���?m�Ѯ����e{l��Vob�UBzy3J4��)n��E��)�x4��ǋ���2�n��n0~�������J[j�t�9C������ �E*�:	N��cj�7�y�pr�P�f�)�UuZ�/+�Q��<�A�� 0��Xs2�Hz[|�1�3����4�\�|�:,{!s��٬9a}ۣ7�`]p����Ǥ�q^غ`�O�䱼�u�}m-#��f|�;̣=$��7��WB���&�n����}��~Tw�=�7���\�+���3�"��>��D��6��၅1�p_��q�Zɲ@�����gG��/i�`j��䦧�Hɨh�4�Gr�B�{:\�9���kl����ݟ�j�&�D���k;uђ�!T^����!(VH�FL�,��:��)�=V�NG[4h=1:�P��`�k�]w+�V��Q�r���l@�S��]�*���į�߄�Xl9g [��wX�h|�@F=�� ���L�����X|�V��M����cQ���;�aɵ��fr�m���m�A�ғo�h[}�F�շXlxVHYEB    1e12     920@G����:���kLa�|���q���՜�O�k�J]9+t��g4�s���D}/��綁8g�w���">�Q��-o�3����9N'6PJ���kw�����l�>��|<�^���&�S�6M���On^��);(0�I%�mV������Rz"n���Ul���U���2�0J���K�c�w��R4��,d�Q:!Y�x�!bt�*,8ƞ��0�������
��]�C4 ù	�G>+����؅�a6�i�ܝE�z��cS��DR�^��Ӏ�=dd例`���r�����]���wX�/����󆖠K���u�;y�W���r5ݤ�
)���- H}��84r��\�
��>��Y�����Eu[b̏�9�L�Xᨌϛs�o���W⋔9WF��i.	��e�k�'��v�aَ���/'i��3�l^����%�B�G�ED��l�a>f��@�A�j����d���G@�A	���O=ƹKޭWg�0�!�*��\�@,k|��x�vT���x�zή;����cbB�lR��"σ:���� �7u
*_�p�9����0_N���l �l	ӞD>�Y}�)��(҆kV��H\7��a����U������h��7u�^ѡ���2��˚�F�z��q>������r��.1#�4葓]��,}ͼhw�cc7;N��XmC�����=�8R�\Խ�3��=�xu�!������Z�L 7Y<�	:�S�� A���A���diG�Qx��Ʃ�1�/��v�6���Si��^��^�d3�5~�O�����C#V���cPc������%��͐�� �l�:��b	mǊ�M�b��^��r��6wt�� v���mJ玮v����[f�g�ߗ���E�׼����c[�)���u����CI��cNd�D��{��������gI�Q�yo
�uoԈ�-�-�1{yq6����o��0�Dj�.{��"񽤰8�{"���s�s�:�,n�/�{��Т&Ym��q�5�M�����7e\\�g�D�a�$�:����h�/{�];y?Bw�ӲՑ/��!�6�p�!6� ���ߪz�F�m��R)8��m�Ǳ��1�Fhm���m"5�4P���vt<$�έ�`m��u�suhB�O�����'�A����9���q��W���dIs��i��8)glϚn�6/=�A%���r��G�BƢN~��}X�������^fSe-ܫ��)x]l� W5P����k��dz�'�UP�*n�䎫����(�s̩���F?O\�픓�Jh�`�*�Mve��1�l��t����9�u������iD:qz�k�na�P���|	?�r����h��8}۾O�������4����u!E�$��2�|�/r��ζ��4��V�f0_Vb�_خ���-5���� Zn�����v�&jȫ6�[>WVv5:��6mI��فڕC�g�Op�6��۟���~�!�<ӷCD��pIN����v�n�să&F�4[�t��$��*�:$AIa\�H���e��;I+N�ԅ�&eІ�>���S�zL�.~]��z���?ok�z�QX(L�ť�Q�?���e�Bpx�����pϠ|	]���}�&��Y;��t�!z��xvo�M���3�~���z��;��
q�~�mш\�5Q�DSz�e�������x�o�;em��ƍEèv�6��5����l��\��\�����|�%՜���,���ȏz@�:e���C`�@I/1Ŵ�S� >㦋�F��)�5�~x����H%�%7��؉�P���'�0J*�B��"��w�<<��U0_Z��k��l��KfxC�)�9gc�b��V!����;��}Q��H�*=eIZ<���1t��s�������u�J]Ư�5��}���4�C�����)�o�2�y/�[�ݜ�tKٽW.� �l�Q��NgA��h�Ї�Ӆ�2�u�4|
)����qp�=�f'��Ē>S�#��a�eg�r�'rǳ�?Ď�?��gVVƣ���~�` 1��s�!fK��jߴ�����f�}��:�r��V��I��;���e�����	�\�m�#��1C]��_uF�Ơ���wI�ZP2?.�[�^��1V����z��<J8X��?��ՙ�掹�9Wվ>4z����b�݃P��9�ƹŌ�ôǁX�S/�g����1��V=�.��Qȴ�ֳ�VY��^��e�m: �<��JC(E����	�2�0S~�o� �!�@������%�� *�j�eend�S�L�e�o�}'���Y��D��^��C��"���7�