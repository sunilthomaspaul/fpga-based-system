XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����|8�SN���h#�I�"M^�.A��K	�<�)����:��u1��K��d	�gЈ�:f[e��
��NH�J;`�ލ�uE(�A��4�-��~0*� ��6�1��W�Ty�:HՕ�B�M4������ʎ ����z�v����+�,�ym�ʻ=��PT�fO��Ж�FF�11������A�U���4����V���YG)+� �� h5%��;�D��� u�o��~����8 �����&����YR"T�n�ީ�&�`i��qgSȜ��ic!�I��Ht�%\^��/tϿ�B�h�ZRG�ĝ9%��)d�����.P��.X/F}�X��W���D|�[�dr���|��I�J��g�yU�#���˶�6T���'͇2��ށ����P�� ��4��<��S�Cw~W�v�Y�+H&������Z��v&{�:r�d��w������ЋD{2��y�)��$�'�;R�2}"rU��D.ўx�1t��2.!��V ��[{��py��9�H.��^�`�`��dF��~>���5po�PwTR'��lT �$�;�3���e����ɳ��h��BZӾ���8F��#1��XMO>i�4A���8!�M�w�b�S�)�� �_�?�)�R�S{;�t�������@��#�%��C��R]K�~kH�u3�{�.2��r�Є:j��NO� 9j0עf��?jI�c`����K��ǂ/�� j`��ؽe��%+l��d�\l���f�\�����E!��&�|��6ռXlxVHYEB    203f     a6078Jy�(�)�s�>\$������Ǜ� �j�T�@]�a�!Y�'/��y��>:k��> �R/0��@�G&}DΕDI]!�M,���������1���]g֤�@ޭ��m�~���c�b��K�惕���2����V�}c,��US�2^f�o��]Q���b����w�>�B�W�E��IA	Ul����-����<��C��:I[�Βp�ԁ�Jc-��Y�������~���Ư+��:�h��Y���S~�E'ev�2�yV��9ԗł�''T��;y��9r0LSO~��7���%����{.7���S��|ֱj�}_o��G��/��΂�L���]M��s,0��~�P���Z=�O�9Cq_��J�PW�d����ue�IA�S؍�$BƝf����\��/!c�j���^��D��Y���ч�<!�4a���I�K9b����8t�b�0�Q5/X�[y���2����l��I���{��J~���$�q �}ik���)�T#���p񢻡(�
�V+���+�'ϔn�S~����>W��y�P����8�0G���[ ���K�4/<@\3G»h	��Z^��:����������.���ꢸ3����j��S@����(�R�������Á� Ǜ���N�0z۴2 =?&�=�Ѡ�W��h�g9���-c)�1�W$�n/Pzت&�t����hN��h��ȡu�ر� ��֙i[�� 9[����nĵ��A�H����)�E1'���!@]+�"d X�;c��Hc�B �����>��C�/�J��)w�������H�s�=.�JTߞ��yol��٣�$n����ĐE���(��?�:�\�a�0���1�6̋��Kz_�\�c�^NN\3 p BZ|�]�jKH�q��l]��,M����ϒ����n�x�'ұ�(G���6>3FD��o)-�?F���	���#<��L&��Q0�C8w�E����[�=CX���7��ц�����°"e�Z���3gn;V��ߖ��^� a�(ލ��bJ�:�"��I�c�/]|i���]E���q;)Ժ�Z&K�F]y�"��z�E��]��@�y��ڞi���n;.�M�I��x��:���veLO4嶉�p�;)�P\{��P�D*�
��z�ZH_Đ2�Ǘ��e�>�jU����;��zZ��rhYyz�?�WP�_��rL��27��]Mx-�	(ltb���akL�kH ���	X����zp%�*�t+-��/�&���|�z��A�7��$�R�
�S�'���~	o0���izs�*2�nڇ��!MR�R��bƉиJu�@��U�9�u��Dr����8s,���]h���")fmP�{�|�<�_����W�`�¢�H��sЎ���{�`_R���H��0M(,t�f��Ys�	w��A����lp���81�WJ�8��*�h+*
�t�ɧ���]�^S:��X���8���F����3�ɤn4�t�^���e���|�K�	#.�Tp���= [rV`��y?!����[��5ys��X��y�����#'�����*eC�V�e\�fX��Ŵ�؊����l�ۉ��_Ԧ��_�9:۔�s�(�b^ܸ*v�JD����y���Z��<����b���'�:΁�֐��V{�	�A	��8���w�K�ou��,����B������R,POf'DMca�ۭ��Ά4DU�������gq����ZO�6S�nX��X���7Y�
���s��UC$Qw$P�L"_E3��bA�QJ���t�_@zxI��Ic��b�щ)��[E	7�tZ�Z�oQj�6i��`B�G0��ʘ�p-v6�%L�4�PKG~~x}9���u�S�����H�0sR�%�-��d_4y�V��r���_8\F'{uGϢ'��F;�Ѱ�9^*�?�(2���*Ϻ����:�~��*
,�@����� ��
���)��� ��xoeOkG!�qnn���O$=±�7�=���MvY��U=���̜E؟]��>U�l���u�(���QI��0��w�]̡2D� ���Q�h�F`#<��:��G�=�%��c�s�J?A�d'� �MA�Z;wW��=�' U���K���ׇ�����P*�Y�פP��2�^ʤUm�i[dC(0�Ҿ�f
`�	'g��	Rݯ	����֛_ۆ7?���T�i�C�v���݆@:�d�j�TvV���;,}D]�>p)�xm�}s�ʃ��p��qP�{�,���[w���e�%#�Bj+.J�z�[Y�.��E���X�L�XhU��X�zv��q�V�!�Z�d�5�� KQ$��1�@D6��>b����٤��-��m���֬�c�SQ�׾�0��쾳O`�Q��笩L�	r`UL+��{r����┩Z����<����(��$'x�a��UE�=��;����W��D+���1f���g*]nK�a�aI��������]˗�eq����Uoa&��t
�q��U�����&�\Ԯ/�g��H<��-Q�.h
E*a�P��]:g�UYt�u���E;\��p�:�3���%ܝ�����Va8c��"3n�#�97c҅�&�#��z5B��J+��}9