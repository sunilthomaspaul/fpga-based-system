XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��F?���&}S�����{��{�f��4�b#��z�t��6��(�r�8�~�M�,*`�	a(g�xߜ�&�lx�G%��d���<	�W�O�ī?��cIT�w���n�2����?l56�Rwo:/�0���8LV�ˏ��1j�Z>IS��*��}dF9�v?��ö�����B_+�u�^��N��.���W�����G��[9�I��2B�;�Ղaa5��"����KT�U��a��d:�W��*	<�4��$P4�8�<� h���n�t?}Ә���'���X,��ɷ-�!!=̗�9��n*]�T{2��@���BXag���7`�z��c>��֥��N_�t"� =�z���k��P�f��9e1�s��O�B�ʯ������
���5$)�{|Z*�m	sr�Ѱ�� Y�_k�����a pU���P�����A�3��� 2˕l��lC��4`�-����'��GC�15�Ǩ��P����A�,VY[�4ߎ���bG�z$xVm�.�������r8D���w�}t�����������1�9�� ��9
�k��Çe�_G�9����a��K�1q��n�U�ㆡ	��̓�E��刧��k=���Z���mO�.e�yr��b��.+������Þ\/  zȔ������g`�}��_k�0Y���=ލ�k���g�8�7�"�d:sv0v�Q��w��2b�����n-Q�U,�1dD���T�t;�74�������m&�XlxVHYEB    3292     b80����q	����;cqMT\�P��QNE$�J%��=_�O���������zN���ġe����6X��+^V�(~�GD��`�{�0��p����,O�A��|1�0�TcLp�V��e4��Bl�$�>�tP����m����g�#kL�M���y��R�R��vk�?x[�y���@P�{�-b!�z�$���Ѵ��̄�xBg�r��~��1���lQ�`���vP��*`f�X�4��SL�]#3�Ypg.��~��3i���Ows2	,�E��.X\���m�U�f�:�e
�diƟ��q�O���硵s�v�r�,\6�����k�ѵ�����T�bW=8��kp��?WK���d��F�Z7�\g|��[�ӫn�&��^�f1e�~��0�	�@�"9��؁�u�&��{� ����h*�ax��	2���̀�.o@pH���M7�C��A`��{9�=E'�S��v��
����b�7�:���ε3+���iL������;��}"�i!!g�ي���2�8�}�nC��{bI�������d�KU!�@}�G���Ӟ�~.]�k�1�����M)�{蝋�J�Ɵ��� m���G���Iubq"b��e}�:wŜ�yob�(��G7�=�.�&�ə
͚�R+����+����.c#lծ���Ñ a5��,�g>�W�K'�X��V�R6�}I!3]y2g|F<�t1�!
`�:��h���/���&b�k���_�f};���L����K�a�vJ���C�����Y��I�Wj��t�+�s�p��&r��gt�K�RD�+Q�a$�8���i�gI>��u�BpV;�qϼOBp��FR
l���1����٣��0n��|���F~�B-W��4@�cT�$޴B�T�P��l^�c��JU5�2'�0��"kr�ȉ���!��1;�+����� �{8��w1�5�c�D�d�4(0�a�eM��� �wl���$t)�ʆw����wB�j쯎Ѯ>�,R�~�"�K#���M��n}Ꮘ2� �̎�lNbs�^fuT|���>����K)X}O_����G����+���[�+�/�)ܦz��"�KM�����p�)�r�u��G;Z哦�E��)�oD+`�J��\˳L���B�W�.�*⵼����Te�������s,����r�s��'�/�A�þ�����ջqi��#��A!I{���|N�6L�#��>`�W������W�>lC�Xco��`�����\2�P�	��ľÒ��C�#�#� )���S��ayUZ�ħ
�v�'��rǽNrC��Dpf c�C`8��=�0br�q�Y�F���-O�kv:B�f��٭���kW
��5_9&s���8�;[���������:�Y̪�4\�ф���I6�_o�9�V����1X�b'sĆ�h�	�iU�������2�ؔ&��v����S+#�s�.�R�\!dnu�[,�-�[��
r�98�Kk<�|Z �d�(Ҩ��R�"Ift,�PҌ|Y[��](�S
�[-k�-�*����� ��Sw▽�0�sv�����Q��q��V'��ug�We�*�m�O�.�Bkx�Wi��pW�}3a �y�ߋ��W$y��=�!���9����,&��p����ܪs7����˶���� ������^Bd'!j��M=Ra���E3����LX����_�h���:ze<��	-.�IQ	I�fS�g����2�� ��X��Oͩ�!�l_��"ͻ2T���ʤ��5$���Jj��P���`��-�|���g7��f���c��"����y�4p�y��N��hӾOș{���J6eK���X��HDR��ϗٯ9�1M����ݚ"PR�0�H5r�����뺹��"���L�Gu�b���9����.ΪA��'��^V�"V*L4��Y�����@�F���|�D�&Mm�9�m�zA�#= g�ٳ��Zi�8d���~_�ĺ���a�x@�r���9C�;<He<�)�v�³�ժ�)����ϳ�oO.��B��};��m뤘��YO�`����O�Ud��	�T��)�F �o��G�8Ɇ$��:A0����]c�x@�<��0r�h��oXҧ�:��d��b�Z;�~���Hb���_�8~q�e;�]�C'����Z5�~o�J/�[��h���n==������p�I#�הL�����Dɮ��4
zՉ79ã�Ig���\�4��r�D����K�p��_,v��^���*��-����%k+^���Q�d
�'�}e?@	�%���k�s!a�)]zM�w��o���qC?-�aq?϶^C��G��?4�}J���C�@E�F��$W#�#(��S�x�R߱fl��������*�ϸ��4'�A�e<�w�A-6i� NV� WGog�E<mB$ �ŋ��?P���tr��P �����Um��Qw��D,�ߝ�
?@�ء��@�#�U9����.�Ռ�H�9cE��.	���������ZRj  Ҕ? �@Z��>����[�/F��A%�9q�͒�B��<
RJ�w��Ď�ǌ U�Եs��"��37�f��
;�*�.�U�eLg��-غ���A��MJ�,����V��a���]Q��e�3���_�D=�'�E�w],-��}���a#�&�ת-�v���wJq�|��3��(t\]]��{������4�|Y��.�N5��"|kH�{E�a�Y��p��Z8`Uli��˵0\9o���mc{���J[l�bKJ�H%��̝�֏� �cK7�sG�q��F�H�L5�c�(���Y@�:T�x-_,w;�؁P��^���
ws]��ӰRa������V~}O���$�]8gwC�;�p����%靓l�E������h����n�+E3