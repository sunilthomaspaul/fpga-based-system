XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���[,mh�ն;�X`�m�6�/���k���سxQ|3�	n�ݛ�����,�=wڻ�ޢy�=m�9_�� �𛚾����!O�5�2j`Ȭ^k��J�����cd���b�ɮ����CSы�
=��K	��3�d���ҧP-\Q����,6�OTMv��CC\0�z���{��.���ELƀ��_8#�4�W�����-g�C֮!xH��U������(�17���H,:3���*�Xכ�#�V��v Sg;���n$9*@�P�Wa�3?�[!�MVn�����q�A,7	�V��hia�t^�7%���ۥs��(���������F���1у:���$B1��ld3���U˒�'��|�V��N��Y�oo�}:;gW��N�q/5�wI$�f����e�^x�aC��Ʒ���W\���G�a�dP�✢Ԯ�
5�j57�b�NmHq�]���Th��ZT������of�<]Bs��K�D�%�(�O���/��D�H�7�2�0�`�7{�^!1p,_�H��*9�W�jA���ae#���zچ�1�A)�֞17������C9v�f�W�����z�WQ�Y���đ�A�iE�)Z�ʽSRteF$	֗ �/RmP�9mv�������3U#�3���5�.�P�GK�,�O��%�qX*�=�S�dT�
�/%������9<�3�urM���[����B"ˇo�oBp����^�y��ϔ?&-���0�4��6f��H�![�� ����::ЊdN��XlxVHYEB    5f5a    1490�Ë�3j�|l��-�8z08Y�=��_Z�ꊷE�п���u�u}��h5�E�c��[�,�$�!a�-1��5�j���K}�1�q[� �#��-�b�Ϻ�A�A�# ϑ��#���yדB�a�jr&T�"��-�;�ń 06X��ީ�äp@IE��\�W��iLT_}�a+zj�q�q��[tH��{�l(u���1*{5Ș�yc�*+�>Z�fhqu!��c�W0߲�{m�`�i�NcT����"]FѶ/W��uL�#�O��׬�հ����(4Oi�zNb&d�z�u_?r�T�g���E̔�N2֥&1j0�xCT��(�6J�?����.���P�a��By��A(.�2s�iI&���08ͣiI����K͖&�!��]�E��|6��^ò1�*l1e���4��;do�G�{��� ����@H����ds�*��~�S:�f��15�)֯�(��U�|V�j@�Z�K�%��JJ �Լ>t�L9^�#7�g�vfL��I,z���,'��n���}<o��G˥�V�[�+4fGU����(�(�V��7�=� �2T�S-y�~��1*�#D����0���-�QY�Tp<��U�g;H8e�Ǻ�� !�ޘ⟇�qָ�`�]�U�����2��0y�g�g	a��j��Ec��$RnN^�2U�4S�^�1ű�9�
��Bx��@��~���n�&��;��9�nc����9O�
��
l0���!�c�Ͱ���>S���k�q�ГV�ru�}݇d5���̊&7�����1.�`�J�S4u���O��*��u� ���>�[|�� �ԖJ&upf�{P��\��R �PG�Md��0�(Я�&��f��z�������Dz��	4htm4�����8_���
�Ne�؋ʹs|Г�bx1"��j��10H���&1da�M&�v=����i��C����/�s#O�1��
��(�n��38��F`��5Bn�z��"U���0c;W�&K���n�܆���R���焊�=�g�uo٣B?{��{���A7جG�d���;U��Aq�B_OY'ZX=lyo�B\�s���9F�@"�A`J�9nL�Ż���w�ԍP
�q��:�h!�L�؛\2�����,��g8�7�S^񲵆���Z�M(z� �.�귢�M%+�S>����N@Z�ޛ�z������b���$�p�(eF�W��%�
\���.6�k���'�bB���G�#�R0F0�E����n�i�e�ښZA�9tW"�52Ϧ�`��xQ���+6y���t
�)i����G$��X����N�6�s���@�IҲ�
���B����#�!#�36{_÷�<Ur���P����Ɣl@��L�Q	����� �be���J�#� �3��H�|=��5�س�W���|-olɲ�v+N��fH��/׾k]-L�:m��u�:[	��ͦ3e�wT.w&d��ߡ,2�;��B��Rn�6�
^��h�@�}��6���<��#yj]�6��ߨpr�z	a'hT��o��%�^��}Ȃ>�����7T�ʜ�C$�]���˜�2C�P۷�j���y�=1cѥ�԰Z���"��POG������2�E�\�k�ם��0 ���� ��A���������<�b�F;�R� #�;��X���6lŅ�~�o3I7dr@�t~m���6���v�� �{1���kx Lr���}]�ChƖX���/
C��fbѺ,��$ݧ5d��O=?�K/�h�����[��Fe!�o��c5���L�͘��?���X��a��&��.~����O�Wғïܟq3�Q^�1�Vs��E��4�
"*����	/.�4��Eme-�J�	��G2jwi����D��&1Ҵ�nAT%٨?�z"ɟ7S+�������DG�� �=*�5}k��.�"�RoF%���z�� ��>-�0��i\:�.�C�j|8�h'O`�ˏ��G�
Eli��
[��eE>����ɑ��LMj��}s%x��K�O�N~���'nq�a����Z�-��4�����H��*
q���]�|.Z6���Ĝ ߧε�ME��9��<�mynE�4�R��vjtZ�`,>Z����)w��?��夑ѻ}�?@�-h>iOȍm�t���cJV/b�]d���|r��g)���m5�zjj�1j�s�+�5xBU�����]RK�պցA	���]&�����z�BW���+c��#�3 �)UGNU��Z��9�9qiT����~�as�?}����4��E=A�w����Z@wD�{D���3�������uL���閭���=9�B3�۫��}|��<�$���(�N��{�e����q��:|h���b�wȶd�TI��� �"�M�G�y����G��.,l���kɟ�.؝9�����X�B-��W2�����3���su&��g6܀��c�P��*ޘ���T��^��j�2\l���"!�|�Y8�Z�������Ҷ����;��_'BY�}pM�,�ה&�󤚂I���48i��_�{_X��c�׵�Ղ�zG�C?�;簟e9�����1�<�e�^nA��G��g�lzb�Q���[�U�Bet�/!��d��p��<^kb���>�Teܮ�X�I~����J�{����N,]���vl�,5G7fe�/�ɫZ��}�(����A��aKȎf)���"�e��A��5}5c\�v��ˆ�%�T8D�ᵩ��h/����(����E�����6��6����� �@�����ה�k�r6�au`̀�M�(P�j�AMoU9��Vb��4j�aӬ��v��'�tM�EU�<`�E�&m{��nH@��Z2�Y��v�˰�����b:��h9݇����ġv�ދ���g�u	�����L�E�?��_7��&��+�Q��`�<�����x���{[ʲ�NK��L��9�Aa|b/���>�c���~���Gz�w���Yt��p�!N��A`o��?_㒶l�ʂ�.ׂ�:'Z��ғr<��yЏ-�A8F���:�'��C��=��0H�3�Z�"f"��{�������tfY��ک{��ܔ��ZI�]�H�RlIn����I$�3q)�ʵ(Ӏ�EM���s��p��)qj>/�����G��eV������K�d�rw�K3p���*$,�ĩ���H݋ͳE6[�Beip�/�$A��S�(ۧF�s�E�	{$;'��^
7k�B���Ƶ&����>޳��)�"�Lh����'p��۹��dp=V*3q�܇b��]�b����8	<�A�r��T��֚q�ͮr����
 V$�y�ڥ�	�����XKr��y��كgF)h���J�)�l��O8A<��ߩ@�� �>f�4l�����ˤ��߻FḞ`����Rᓧ����(O`�Um��)Q�H��}��Ht<N1�#y��Y��1�����M��L-����x�ُ��T`t����5`��~����A�>-l�G26�	_�8�s��F��d�Zg��ea����j���(���7h���#��+�07����T���Ek����Uj���a3���V��0���^ma�4�}����OX��C`2G7�꫌!�|Hh�t��mi���ƍ��Fc�9�ܾ��(-�Q)��G����E߬Fq4Y�$�������z@���@kڜ���	Z��! H�B�	aj{��7��d�)@V������\j!#��R8G����幁��t���i���A6Ot��k��IG�_�̧UW���Z�)-@*�We"�y��?��eU��6�+��Y�P*�Mp瘑V�0PU�y��1����%��Z�G� �S �8�8���)��'k���Z_-��H_�:�>G�R|����� ��zt/����w(+:r��_2EU�5Ϧ�46tk���F�r�B0��[r
��'��d�S�c[��l79���zz�x����~2�-�YÆ&��M]	!���c�&��{�F#�%d���������[M�Z?����=E*wG�k�3�x 6t���p4}�&�D���{�����ӽm{#�j��C|���MgLyg=������h���Y �O��8i���R.��@~V9Oaj��A�&CDg����0#��M؎�֖�*�4�Ҙ$��=]����=Gs�I u'v~9���T[{���S���u�/�rز��@�/�ISl4\�ƽ��3Y����:��2���|�}8:US�S���ӏ�A�G�y�b �wX�S/ytw\���'1���C�cy�f--� ��9�6����I��j&� ?;����Jť��Vͺ�R=_�MoqU��� ��a� �u���;�̟S�@�@�ct��&��CڇM�%!�(����%Ȅ��̳�����b�|��ͪ��b5�v���׌�~^#����E�E���j��,�6>��g&?閦(��l`�N\�� ���q3`�S���eE-�=�! )�NC>h9C�J;�H��k*Pc��4#�׫����&I{���D`;���hڛ��կD\ިI{�_��[�o����r���=�����۵��y�e9�/��Q��Hȡ��[�PL��rs���y�����ݳ���g�&�i��^!9l��17&^�=о}��q0G%Q��s�n�[�SB��Ys�&?�Z�f�����f�a� K3���5��G>�)M��8\��K�B��|춌����Z&d|y;͙RD�E*7~��+�Φt!
}d�Ӫ%�.�����z"�,٨�����E��HwH)�ޱ���H^�HM"����0���[!����*"m����Ie6kiS��d4.��� )�p;~Z ���'����٘Mَ����]3��«�N�Sj_��;'�\�
��7Ojk?�\�^^J�n�VulX0Ӫ��G���2�����t$7@C���z��#Ԇ���!��G��)1�eŸmr�@��m����@�S1��ʷ���H����Ю�n�H :�x�7��/w	#HbaG�K}�����K;�p�9�-@f�˚��9�B+`�/��iǖ��(s��o���~�B�)в�F�R\�3��iF�:O��r��3��Gj��x���/i�X��?��A:2/&��ۭKE�t��:	.�E܀�;caL�w���j�$E�{J	�	ߜ