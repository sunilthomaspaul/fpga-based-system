XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��.
�?fz��{{�NP8��<���Z�s�hL� ���͕`ߖv��T'�S?��.�"��p1t
�->���B�m���B�ñ�lv3�-NH��!�
9@��8E����ȷ�V�s�6�q�,����d*y�ڿ&���/p�~1���e�A�@��O�G��7 `��Ѥꪊ��B�/#�c0xKXnt�Z�q��ó�̞YM�z���x3n�=���vGF?���"�fn����w���O�^���	���q����l^�J�����L�FtL��Ҥ8b	Xu窞N�B��/	��G*��6�����5����o/埇��9�&T�Bǆ�=��'x��j�U�֙�G=�m�]��Bw0s�]{�LL�4 ������3��EрY��x��$��θ�w�����vK�R<Z���ZRK�NɚXHL���U�B�y$ȹ��[�����n�NnX��Z�x(�.���4B���q����#���/Ձ~w�ceY#��R�^��|��t�����Z;|h��44�\�E�8s�N�%��ϻ�[��"�$`xɭX�/>�F��&魰AP�N�kq������45��o܋������(oPPJ�͇�wS�)��	�B�T���1d��H��r#�{{�5�;�*��2^�d�u/"U��c�|$�<K�xa��C4wzY����:�-1�ƫ����n�NR���� b��(fşm���=���j�!8������T�͵e���2�c��!������m���XlxVHYEB    1017     680�m��Ѽ���]�mG�0v�YA|͛Wt2�a�Ig%W�l\>��PFh&�>�j��/�;����4� ܑS�д�v�Y���4^N)k�CB�j	��lL��$��p��Tn�V�!)�>4�Cs9����K`�PW!�����8�����kr�K\(�F�K*��С
q�����f,~;*X�ܻ{`3?��>�2n���,ʥ��v���r�)�h�W8 e'��������Ț�uc?�qAR�+���ٝ��p�\1$���2q�d����M�D9G���64�e{� ~�'R��r̀�����ޝ��gV�����/�e�3��y���s��T4*TL�ᶭfkCM:T�~u�e="�A���@6�
�)�(E�>�X���u5�ű����>8���A��m�$Qƹj���љ,D�<���(�snf�_;-����.�jS�f���E�kA �Rb�ǴU���KU��=��˂A�w�d���ܲ�cȤ�۬&�"�f��[�ߒzz3��'R��<_�J��q��4ha{����S�F&��j����I[��d1�v�̾��)��]S��F���.[K8+k��H�������԰	��Z ��p����jf��������7�H��BI6��C��,-4�7�e��m5X6q�T�~��K�-�M}�S*�l�ƿe&� ��1�E�����"�o� h���� �j�d)F�0��v����Ea����~;
:$�`�d��f�yh�]�a��]T�"����>J�"֦��oq����dTw8��7᫆O3�츪���|2V	kxJx����U��n��ʔ\[�,ctLu���
�b�͡�6�����	O?���qC�I��~dV�!�1�+.�`4�%��lY6��^i����p<�3��H���<�,���x,� <ka��T��R�ɓsGI�SN�krdx�+X��+n�8���./�!�H
�: FD�-ʁ<�Ľq<�4h�re���!M���<:^���:cP�:����uY��ˌ����Cq`U�?�eXC5����n��<m��?�!T�O9m�;�B��<��п���h�G&�q
�Uk��+�\�U�Љ~̮�q޻�3��7�'�zv:�dM�F�URB�����m$�Efo�h-���&e���)� m�6+��vˆ��{])�[�Ĵ���lSgܞ��/Zc*���~�ޔ��*E�5�>�-0y�w�'wl�4X���T׎�|t`y�"]Z��'��i��W~j2Y��o�#`��S���
�s3��sꪸ���.K��<3�'������Zy�v���TP���R�P-�/(4����'�:+���#��瞲G['�d�C>�l��Sy��q��>��Ǳ��!@x���x��bz��7B�����i�78/H8��q�x��D<����B�1�9>)Nsu�c]@�Ȕ\�%W��4���֭��&�a�!2\7���`z�E�o�R4Nn6���������l�շg����&�����l��Y��oJ�;��\��	@�`�m��Iб�+°� Mߨ�gI9}�9b'ϘR�Yn�B�t���*4�����(D��{s�$�l�o�]�M%�A0��f