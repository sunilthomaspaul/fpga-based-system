XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��@��\>�N`0Y
]�VL�ǹ
�J���W���:��+>��9;���"��ZƼ"��I5y�Tio��ˍ���!��T��*Њ�ӚE)����R�EaY�l4�]�c-KF"D.RI9�W���L����i��CħeR��K�M����j���t�%+�F�E���Ã��p���0�u����P+W�I�b1!�s6��&��q��(�|A������0�d�� �9�.o� 9e��!�z}6<�������!��SW-���&�=?����Y�6@d3E����]
y>���'e7����|��1���k|��|F'-fnP0�[e�@���8��\���?w�w�Ӎ��]y�Ё8���*�����H�a�d�1�	*��Q���B&]�]�$-�*vb����ت�7*�B������-/�IwdG����w�d䕨I'6�{@?�J�Z=Q���C'�]�R*Y�s���/"��ɨ�f}��;k�ڎ{�l�b\��Y�$C��=�AlLoY����JZ����w���R���:愀w%�p	���dl]��N��J�`[�t�����7d���rr>�9._�����7[ө~�}�4��J��J�
���~�8mt�|Y8���#��6�t�g��A���΃��V��#vX����m(%�AMGL�Vى��y=���l!�Kjd���]��vU��(b�09^�_R��E�|����c9\ģQ�|G}eQ>���PG��s:$��  K�i�XlxVHYEB    6ff5    1760G���i"��!���]�R�^Q6�����\YY��u��u��O�J��~���kG�=Z�f��:����b�4�m��\CA,E��^N���|�v6/�4x�Ƶ��zCW���ۛ�&����V�'�d�	��U�&���i����R7B�y�O	�w�疨�Y,d�k�
$�V�ݙ90nX �cYAQ���^"����c��
.r\�ɘ�u��1�q���7J�vrp�[-%���C䒇ED���<v\%Pd�T]c{-�~_�R��EB˓� q�RَDh��Q쯹.�&����1�O�
�� J�pArr�޳����KpCr�h�8��m��}�������B*\g/O�v���k�;���� ��i��X�{��6��^��p�Bv�nʺ�=�<�Q޴�]��q0����!t
~=���b���&����X��ܪRݿ�nǾ�y����1M�9�F9�#���M"W�`2Zr��e�"��j���,�^"��E/�y���1�M>	�
�<�=]���> ����� �C(�2GT<�����p�\��AyR,{��J��`�^�,����wjf{�x��zGdy�Ck��W�Y�xFxt�R������w��n��������V;�7�Hx�LzY� b+����ͻ��`$���U��T�)e�X�ͅ\�V�3VX�A;�q�&��)R��W��
,���Y����[+�[�y�7f��bܜ'g�?��_R��֐���e����LR�I������k�����1�{��U�\}�_þC�u��8��2�[��z���S^M��|b2�6W���Od�,�:W�'n��|���!�J���G�<\�0��]6@׭=7��"�?c���4�6��Jb��ᓉ�v�#+Z4le]|���yڊm�!���7knD�d�y4�s�L�}*8Ư!��o�� �v�����i���
hv4�z}[��7+�x�BӒ�(��,�<�}��yb���������i:����o�nP^�	����3�2�0�������(���*���~�2A)_�l�R�E�vX��|��L��r�<��~��K��U�8���<� 31L��(Wc��SCͤu
��j0���T���j[l�����l|��M����PD�`����}�~���{d�:��(���LtT���f(Jt�8U�,D}q@{����x��w��%�X��8Xk}���ꡠӍ��7�T��C�g�^��q8b:� a�u|�B�� ��3��sC�]2�~ڬ�� h�cjB�~�8w����r7򩩠�~�Ôo��g��y���q����A� s��~rcϢ��V}��!�<�30��ay��<���4J�t�b68���)��3`H�Zs�a`�s�E�Њ����T�W���M6�l����c;��d��S5ߞ9�V�v?Z�H_����:I�-�_ƃ�RC�n�I?�UW�E����;�6��ܾǉ*��a/J�,�l�$��h���=��%y�JgC��;�ժ�)�n�7V����1��\�6+���7w��&1ѕ�$�k�Ӡ$n_��u���CtR�]�*,�ˎ��	NE�ӟ����av�,��a~���n�z3�Q�����ŁҮʸ� ��4�8��J)`beh±&"�.�g���=}���3�1TUb/����	�ia&�xCvt�/��
V9��T�Tg�ᐓƘs�
��D���T�pc��s�����Rp�2���#�)�n�F@�J���:���/A;'K�u�`tpP�Cv:i�B�{a�d��䧷��8��^h%���`�Zy��_>����{q��JE��|Z�x0A�k�_x�_'ǒ\��|8%aBR(����oҜ�G�/�-��؆���*NҬsO�BD��K(�okT�"jXt������=n���Nk��w���3��&O���+�lU���?�'���o.�E��)B�;�PP� y��b��3j���Z��t�9������A������V����e�?��+qI
�@T�͐����7ng8�z}���{�~o�)6��5c]�]z�-A��J?��iM��=��()�r��չk��|AuXM����O�%��u���p^�}}(5�@PV��տ��\�F��ů1���Z�β��@�m��F�X�BJ�l��!`�_�L�\���ˮ%�똨�0����}�7J��`l<�9x���[�V�(�ї�Ux�f����v~�g��n]�xفq;���w���Ϭ�˽�u����ci M�5q�6��~?_�z��pN�=ɥ�����jT���C��%4��+��K�$;E�a�����*����,�[�w?7�'J��\���� �cL�K��6�d3��y;�eu����#��7]�ϔk�adq�#����4����$]m�ID������� :��^�_��rJ{�#��������:������YH�����,�u�4���O �pDm߯�B�8G0k� /V����tn�}W���#�ɝ���$�t0L�Vz^k��G���8��v������$�C �m��]�F��=Q�u6�(�Ͼ>a��1!��I�����Z��|�0�G`�l��I����P�4�OP\}�~�h4���R'��i"�U��[;C�Xӵ�6g�bC_�^���yEwĪ�ع�ח��o�s����gP
�)�:��E�G�ҍgm[7�Ƨ�p �;=��]����>��*)����)��%+�eP��g���	�?�[DGJ�q��Hd͊��b3�5��Q:?�pp���s��8��zk	��LC���>/CC��+D]l��� �SO�B ����G��v�Y����t4L�Lp�:Bb�J��@�kf~Rt�܄pf���x�UZ����s�o��������E8��$����O�&ŉ��_u =�R:6l����G�	D�x���`6�������5a�P�{M���c��n;gW���4�������E��M��e���,�������� ���ȶ�¢؈�z0
��<��>v��h�U��w&e0E�x�-~]�hH]yQ�K%tu�7c"�2P���Xr0J�G�̏p�����3����e�!�����:Z@b�<n�N�s\�=��1cgdѐM��Byv�9��j̫Z�Y��;$3��W1��מ�MIiǛ�AR��aw×���(�yBB���v�����h�\/**I&w���V`�v��4y�֋����2k�_Az��}�e+����ĺO,����)���a��ıD�ڶ ���H��.���D�Va�ό���p��_}�#q�Nh��g[�J�p�K������p
Ь����3�a\�0�1�d�j��5��LR�}꯽	Dj��n�XX]��W��0��K��)�[X\��k�ߨfm���m~�F���g8ȳG�L�A���!t"������_3[2L���X��'U��;��`3<x���9���s]QTY���O_�B¡�$?�'����C�!��:�"��S�fid���L5�ڵ;����G��&��пի'*M�҈�z�(d!	Z��D$�D�/ژ��a��\�ģ��I"��͟�n��=l�9A?Jx�q5�2S��x�ˑ#��e��-��-�s)�
 ?V!iT�]���ԫ5j���Ѷ11�} ��n�a����� L����vG�)=%#L����[kkb��|��0�U$6��p��o����]�S2 #-����;d�"K��f�ub�Ja*��:�"�=�pz�c�Oת��u˥ɉr2	/M.�6�_k7�g7c��Q�*�Ը������ �O[`g�1�=�(b���?�}�@��aSc���̑I��@H������yZ�)���Xf�4�.z�8A�M�W^��!�V�@������KU=��Boc�Ƿ$)�_�nd�=e3��i�1�f�G��,��ɕz����"��
+EjI�{Cy\��x5.���i�哙t��J]_���qJP��v�Zo��d�6/8˃ܩ�u�ϥ(�V�R�#�;yޱ_��O	a���&�/�i!7��'8#?ӿ�����ٗ�@\'�8 E����`��?
N�*7��̄-�������$�ו:����V�$��!]j��ņA��&��L��%�O��㎊�6�ɜS�b���ɰ��8�dؙ�Ũ�p0+Y�F�;e���c?�[��)1�L��WKf�=X���^o��z=�TߛɜR�0�ܩP��`���?�9�~Mà\j��S�۟j�]�X�vZ�?�D�4\����|�S���4_���T��e+K4��{B��K�by��:����U����9VB7�:�x_'���WJ���"F�"h�P�jG(�]����:2t���v��wDޝ�=�B�z��4[Ѫ��]���]#���8�-��){�0�=Zn��~썖F��_�)̛�b��߬�qpU�Ba+?2� �>�WK�p���7��.��Ls,FN�b��K@��L�z��A����p�D*�Cۻ%�[��^���PZ</ǩ�6`j����\�H��?����R.28�F����1�߼�3Z���F?�[���)C��0-&�j{�L�3�$����O~z�g<�s&O��<~R�>rum��)� t�@xĞ����M\8�7kN,}"�*�╋Y�Ee;+U������ph��
We^8�,{i�Љ� ��+�f~�^tp������ �Ό[�>�d-%�]L����Q/z�3}φ�9�RL�
���f�߳ݖX�z,�{R,���i=�N��-8<�����7�� ��2�B��c��6��B����5Y|��6�J��T�
�	��'�O�#	;҈AY\��Zv4���_)g��cxvx����;I`�)^�v�0��>)��>����;'H^/�-Z�Dgc�.W��3ܞ���B���<F���*����\.��+�5���k}x�.V3#�T>��?�eO�?%%=��+&z�n��*�ݼ��&h���S$βmA��6�N���j�xh\5��&
Q��1�H����I��)�u�Q\���v��F����E�2g'I6��	Y��4�]����c�u��XK�=�S[`}��:�|97�'L���k�2	�c�y��� ��+Y7�D�@r�	Q�,�F���$������Aw���¹W�#jYY��ѽ� A�"�1>:.�2��t����AP�X�|�񡘃������<����%�*�M{h��� �+ã�yH�k�l*�26�f�)�:�jhp���Z��C����H�K:�*��`8>�F��|�6B��wߟ�]��m�+�+U49 ]���S����E����70/�^k��� ݜ��53���&�'=��p�˚z�H,"��h�8@atFR��8m#���ɯ2w+�i�b�戩KgC�a+�n,�����A�$�'(�5(?!\�tPp��^Ċ�j(:-{:�d?g6�9���7�t(7%�}�q*�?.4xqJFq� �~��>R��nbUI��c��T)qX���I�td��N���4����wig,�F�9���f�:�$Z/�$������y����?8B����tձ��RC��]�Cp�}�|K	���8RP����/���y[r����As�ЧQ�J�M��>�U���R�>(�ح���g�����e���w��ᯨ�R�r�Y�Y����*4����'S� �p��ߝ_��V�n��m���"��1��^?kI�dԗw��\���g2��;���Sg�JP��:?e�ݨ��G�C�J)V)X�)��>�������wݮ�?�	=:���'��V���qq���	R�j�q1��q�d�;���헬�l�I�#��%