XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���l��Y|�B���7��
C��NtM�4��2���Q�����!X�I�Q̯J��T�b�c���z�c)�,� �[�#?[�Z!��A�غsk��4,� G2M�{�#~�xn�������%�+����I3(+�{,��i@8�KҞ;��.|}����w����0�J(�����/�s򆨃��,!)��9�+�UĮ�.�l��(���S����ޫ&y�����PXnqi�=��*N
�$q1�)�����'Z��U�9�&��ǁ|��X�
Ȓ�&�z��R`��6��	��Cv�V� Bq���gğs�u�4�㑉�63Q��]EY��y�.�� ��;����G�����A�KN���l�+7�Vp�83ɝ�~vC�=���B8S7�KP �[E���<���f����@����#�7��~su��)����������Gl�l�k�zb*�і���_��꡴,��<��dÃќdY/�r�+P�ԬW���LWŧA��#��8�s����@��|���H�~"��+}%�G�%������ |wHN���O�!B�����H��i\����f��\�2#�I�!�S���|��qj"W�J��K~��S|[��}��O�,�1�������]*����ٟ��W��\������-9���S�&`H�G}"eJ��MX��OCcJ �#	�fv5�-�tq��wIBBZ샎��t`܅*����r�+��W�R��Wk�0�^���q�o��Z���p�1�F5�XlxVHYEB    5658    14e0�1S���w���g���,M�6}h�_n<퀺N��,@�^ c��[N�k�՘|2k�?�2�$������n&��<�m�垤-�F�v��P<��8����(��b�π�֯Ӣr�k�?u'W��b�N=6��\w�keqx�������̛�/��1��9�@+B�v ��������?�Mb~�������� w�>�+Q>T���	n]=y��	=��N�o��f��Ah9�w��lN"�����ak/�טʟ�Շ��ٲ*\����g6	ʢ(F��&�/0�:w3]g�z�Mu��uqG��8�����H����0p\K�Bt��厤F� E�[��{w����7#�8]>$�(��u�'�w$"�a�C��Dd�ວO)-�s�����R"b��I6u%c��i�%+	�}���Q�wӘx��rSk�4�g�"�u��S��m'Zn�/�;���wH��8#�8��̲��e�������M��N���UR��v�\UUى䍍�d�OAb������Ty/�b�������Ywt��a�ѳ\&w����� X��!(|���؄��_���l������a,t�l�7���%��� �u�f�k�����9��1�o�cA�~�EH����}ےF��?���r,�R �f���� E��o��U�#f�T����-��ߦz՗�|�'W��s��(���A�;.�W�yF�h��������~
����R�t>�7�k N���GlB�����U�_���Y[ྀOb�$��z{Gyl�L�4�עˊ_vR�����٨�񚿿s�X;��3*�js�c����V$ˇ��v|o�|P#���J{h}J�C��[j��6ebF��u ��<W��.��u:NΦ3_5e���e0G YZ�mE4�Tm��F�*�f��k5��(�;�'�b��҃UW�?7��-�W��ć��@�b�汝��|���q���v�N��^>��@�T!f9���-^I!6�URN����lJR���V����&�l^���ޱ��~	-�Hw&/|��B%7���'��U]ܢ�"����������b����̖,��W�A���xTf�(h��@h����_ʶ����G�J�4��.6��p�#��?+[C�p��ɥF��z��g��XGY�*��v��T��C��+F©�}��a�*�k�/�X[�|���a�јh`r�)�����R���:Ũ{�f���Dnrc��4��n�/0?�V���%A�)O]:M�̼�F8;~��1�
=�C��ꆚ����a�u䍷|ޚѿ��N��&+��Ě7g��pP{k� �SK���:����:M���x�_{{�*G�m��T�/x	�`�y���N���u�n�����=�|��7��<����t��W�~����)S�!��~%�c}�έ�-�Y�Y#%^ی|�/6�u3�1٨�^m
��T�5�K��4�R\�~�d���N�3������gr4Ӈ����"����B��Y��0�D���y�cK!iX�e2ְ�ʉ�TVu������D	x��jݾ��d�=�*ܒ� +G�X+�L��& �%K��5H����-��D�@���r�v�R������7/^���JkDzv'��ʃZ=gO���s� "���KZ��٩F�������rV��#�_rK߸��)�TZ�C�z�������T����R��euda�lW��3���<�/�7�ŗ����b:p �� X/�/�1���Wꂊ�F47�����.?�c��mH���D-ׁ��{2��;Y�-���+�B菹Al6�Z|�Ǜ��:rM�����S���4JEЅ����:�he�h-p��D��7�B�
AGv�P�[�dl��s�i��,�x���uQ�S�)��-�e���+��Ӝ{���>�����:���.�彠7�j�W�y6�ȭx��H���� �x�KFj�D�ۆ&U��३=�Ru�	��l�س�Q2�ĿGY���A9�-��F����븮�#���|r�;+���:����9R�Q9Qk�-oD��Q����s&-�Ĳ�%�s�R��1��Uz��|W��k�E��mc�s�<�"�ѕ�~��'���$����rL���8~޿[��A���5�*��Rq���������Z3�?"B�&(Ni��D�j���Yf˪|Amm+��[�e'������Jn��wq�xp��h�P�� 7�4�1����g���s'���Z%��4�I��P�Ƚ�:�[��E�E��jIo!� B�y�)cz�ߑ*ɂ�#�rB��]�Cg4��va���.���Z������u@�"���+0a0X���׈����_S�8:�gD��w�΢}f_��n��itS�O "ej���T�[���fH������gm���2feˡC��߾��ĮS������sW��?�Ԅ��ج�˾������e�0�*S|���sjM����!_p��P��FK��K%�����v�N�vNni�bFtXW�H)ѿ�ҘĀj�*��ȹ�f�Ď���Q�!>ep���90~2bm���8G���P-0n�7��:Y�_�H'̂�F��b�k�	�ߛ�ch(�>�.
�����b��'X�(�E_`���@-�QV�nd-�L�t�Gi��9�z)Ov�mC���>������K�_��s�4T���YpS?�e���3��E��� ��J��|��L������?8D��*��h$�9)j�Q�b�������d7�kRj-]=	~�gq�L7�C@��6�0����p1ҫ;��zq�Nh���|��^f����R��g앆E�����$�n
�e�����P> e�7����-�<� ���������N'+��Ȧ�Iy��� w�!����'�7��n�iz,Fo�x��?M$T�<��ϰ���s�~�hi]wY�B�&�u�S��#�O�����5 tWUVD5��9zT��=�zJ��3
�QOK(��mi�/x��u������LI�~<%m�K��+�] |���C�.�E�^�oߍ�$�����%x$NC�+{�TZC�~��D��]�g���*4����"��y|.�L�j�b��R���N��5`��~!���A]^�\no=���.;˱(Ph�v�:7��ၾ2��H1V\+0>��̴�Lڈ�9�Z�/��n)����j'2��Y~��2%��6�3k�,���h�0H1��!(c�\իי�ɑ���pG1�+���G7P6�)�P;bE �_EF���v�P��b"�h�)�l�Cb�a+u]6�B�쏘���H�,����h�"C�"'��/��Q��7֑� �����	��$9y�Oa�  ���a�J��m���y*F�'Y��7�^K�=�9?-�`�>o�n�Oz4C�r�a���o�h�	f��I�����0�$�(���z��͛3o�����o&Q֣?�c����n�ak��Z�bIFhl���H���5r�M䰙4L���\
�0�%�TY�j�߻BG4��=���۶^E[]{*�{�R��Ai�PsnQ�|}k�v1�(	sKݠin�ؓ�<2W����%�"I�N)�ͶK�r<�����cċ!>#�<=H.=ꈭ�)e�Җa�Gsb�db+.��41�:����̷�E���~��1R�}�׽و����\�NQ�Aq�<ϣf/Tb[@�9�'���&Z+��ZDU�I=*F������߬�~����?6�r���2��_$�ԋ�?��^�/΅j�,�؅�+���C�EÝ������{p�n+3��Ew��ө��M��RM�J^)ֶ�ܤXHX�s����8*lj�4*������/F�t�"kg�B�8�{RG+�:F�^ir��|��e�ە�"���	�7���+'"��";�k:�#ڀ)ÃP.r���qF_x�O�����	�����c�<y$4���<��>�1�����}��;��G�C0�A)nn;��w��� ���P�Y�)����!����<�l����H�θ,VCz2hF���0��"7�
��)m��]��W���$X��C�\߱A�������t1�}��j���bN����Õ�[v�FђX]�h��z����r�t����|o�0E�������v_�/5lwo�W�U]�q��f"ͯ�n2��|^o�_��x_���\��H&����I�"�l�"{CA[>�c�SM[_K���M�ڱ��������"�v1#�q�91�h&�	���e�`��y�i�Fr��C��U,��(����H���V��@����ch
��61�9���`Y�6�-�%�d̂�����r�i�����W!Y��pS ���2�]�}@��i.pL+ɋ�3�{�֔Sl�L�N�O�X�僫�.>Ƭ*����ޘ�Vr�x��.�a��C>�������O,Z�j�e5�t��%Y�,����6��u���ȇ$���1��y�7�m$�v�9P*����*��2�I�fIw���7tC��&���j�"�\������H�\éM�4�g=~Y�E�u>b�u|n�¹�U�����.v̤͐U���?9�~��Ȑl�{��|�N�8���4)AM��]�8��h#0`R�`�v��2�at��U�]!1�h���Tq`���4����~T@��eB�&a���*�5X���<�.�Ԏ�w���el��l@"��m;@o����`�'|���>)_�+,:�����N�g�g-{!�,�� �M������*��Af*�K8^���85�B��+����ʀs�@ZL�҉�ä_@V�.Q}1��`�
��hm}�=�3k����=�s��w���]�������sur�q$�!����{���tw�����^mb ��֣xP1�L����6����]��'+z~*��D#<3b��y�Y����T���P������k�I\�:�Ok�O��䔨ipbc�nؼ�����$Wu�ŷc]���Ri�·HtU�}�M�:�-׫���;��p���xgٻ6�{L� �m�^���+u`H����:T~\�[oc,g� 2G����7&�������C��r�N�ֶa�I�*U�>}�~)��3��m���+�x?������@)LZ0=g�-�(1��.&U�,eykolt(�l��1��]�$�CKΈT����B2~ N�)N�~��x8��Đ���XW