XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Z��"/KϡC�N��K��!;�&�:����l�Ӻ��	�����X	���F���%~D$�ܯ���{��4wӉ�}Kô�U���ކ]����OAj��Y-f!Y8đ�[2h�w�z�
�@�-�Y���6��g>��AZ��V1XKH�$٦�]�Ip9[[���U*�j;u4�S�[4?u�����m���'��n��%Th4�e-s<�v�R�&f��b�}������E�:	)}ź�L;zy8v����fˋ�q��{Am��]S$�.�#��Q=�]��h[��d���������.��Y�5��r��Y���V[]@�����<.]��u����ם��l�/hM����~I�5N>+`_[�ɵ�7�c���u+#B�ӀC曇@4�N[�[��/bD&�X�qO���wv�s��K�[�1���{�2���(��uR��I"��-�� �^��n�X�2Qv��{(�y�w�����0�=)���u:���/ma�������^:a�I����1s<���R'����U:��hE־�����^?�[y�H/C�3Z���r�N�a+c�Q?*l��o��Y5������*Lc#�iZ��xW\���;�2�g��蜾����/qax�햻���Yx ��q*�Tt�4å���^��i H�?�.^t�GYA�Rhͬ�8ϼc,&�V�ɦ-19�͏�
��%�9�:C��0�p�!'�Lr�{$@Zd��1�X�f���>%����1S�ar�j��e�oC���gi[�_XlxVHYEB     f8b     650���B���.e���=��@%�ǜ�ǲV��(��pR�3bh��8g|~���0 �7�O
j�H����Kp�1��`���������d�n1!J��Q�ظ��\g����ڥ&��uCk��VA/�C��OC7$B�3�N���4�Md&Q_2��[�Z�}�����R^�����Ӊ�t��������H�e�Ӓ��a����<���l� �(+�  @{y"6=��O��6�[ZZ��W��d��pg:�I���/�g���C�8}��Dk3�Md�s�L�ԇ���tj
�3������F/*�lb���|�3�02�0F.մ��:�c\��f&���.'z�W8��<ݺ�7�ь�m�:���<��|w�ch'z>�ǫ9�^q��Z�����&�|YlC��T=������Wz�Vf�	�O ��Af��n7ce�62P���P�:�R�I�iEG\�n��k�����p}|e>+$��<'����>���rw6DbF�36�5\�C ��ك����6B�dl�GY}�wޘ����\#��\��hw�z?�����{p"�`�v�l��>�I
b(�Ud(2>}/3��A_rTLF�n�H��K��18�wP"�c���5��y1���^�b���ǲ�G���dP[��z%R�"{~ƿ������(�p��L; �lF�p���}�zƥ[\tI��u�"����w�i���I��U�z��e g+�U�[��E<�L�
�ʓ�א����$��:I�v���H��%�׵��[ GO3+��n�q'��E��NDc��6�l��?���5��D~��BEtn�Q��SQ��Q��������+�Ȕ�2.-�`�&�?��Y�z$*�^M��52|[/lN(�s����O�p�AR���:e ��#�zQ]Y���10��Lh�w�����E�� {�J�y"ӑ&��)Y�U��G�0�����I��p�
P��`2(�َ�.Z6��߁"���s(W�c���?�!����L;2u���/@$�??���Cȋ;#M[k������_h7;۱�eh]b�����#�#���a����v�$��2O��M�tIu���!E�O.�� ���x�0/���dz�c7��]�&x���X��?ڟ�9�(&��ۣ& �Td҈1�H:�\��y���Q�i��Pg�����V��:�X�>F�%)'�}�Ig���EI�x�Nf$�p�XJNG̞I8�L)�ЦW;��0��.xά(��a8��1�E�Z���("��r�%��	�u)�kg̲�յ�R����6�n8��� 2�L��m���Q�>x»{�ǋ��y�iר�|��Nν��O���"��\c�J��ӳ� �^_�������tnf-zs���'����6#���z��J؄���k4 �9	��nU��(fF���|����/ ��a���P�X��Q8⽍Q�t5�r�@�c�e���Rh���i�%�=iZw(<�>�e.x��^�3����wr�ସ�������H.�YDk�FK�t�f��<�MZ��$4��x��P:@�o"����P<�3}bP{6�Ff9���#Xw�$��s%lp"���ןKG�_�I�������