XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���s9�>��FmV��#3��NB�����y#Θ��&$�%q�G栿�7�yp��7�������c)���.����s���v�ؘQg;j�.5�&�K��$QgI+@�J�"kkR|G#����vh>1��N�'kQ�hg�ej� _S���:2�2�.�=���vP��
��7�镧����()���/���TC.��t�Y�����=�����]���DSNǽvn�Ȇ����~x�ݗ/��=q��KM��T�\)U�FZ��X�rb�r�#��L���$;����Tb1q�����e�J~�S�=ƬS0��Z���Hs[�[��"@i�(ڧl�n����^N���m��ki����Fz[�c�`�7��y AN��
9S��1lO�9��Jc�8�U}!e�Yl�_�Q�ʋ���:��?�+$a�PH��!M���&{YE�Y�1����/�=6{#(gWnf��#�V�9�(��2|�yf�q�V�x�1����v1��M�߬k���|�{�qRR�:��Ք/Ҧ��'��*ul�N>��w�Ң�sm�������M��a�p���*5�Տ`�9�������E����u(8�]�����A�7]��Ǩ���9N�vs����r���`�d?�ao��p�`�� �~�K�˸��uL׶	Nw�X7C2{[����R-�ӛ�c:I�}Di�DWҷ� %�����<����"�k�/l�9�����'���"a��7^����Fܐ򢸀o�kyM��z�]�O�EXlxVHYEB    1eda     880����A���c�]��< �!5�D06J6�8Էi���u�+᳑�U��+`�\�؏.2)y-�T�)�#����_"����=C�t�t$��,]�e�R��y�s��
�g�V�D0��\�yT
���{#3��rs���s�S�H�NċIE
�|�s3��Q�Ƣ�Q2k%�f���_���\�u��HV�:G�t�s�S����[�{6k�T|��a���35�������������:�M�����NhO�~֌3�I�� `}qO&��o��7��NYb���R]���`;b��5�?����ٹ&�D�7�pI�Ȓ�C�)�V�'���ܭ�Ԩ��.�$ ��4������vM�T%��Ŵ*;�ς�Ó������3���|���W�<�C;���5��J2���*��}�0`���A%%z��^<%��0��*2K϶��9��V!q�:�&t�*L~Alt��"3���	�V2���z��-?F��mۃ!O�PҠ��I\\��M�Z�?c3�[.�o�Bu5
��ɵ��Є�N���b
�"?F��p{(�6Ĥ�RȀ��-��gm}�
`m���^[p>�eX;}�v6������"�[;���&vQ+F?��Љ�KP{!�[H�g�]�]D��Ŧ��_�*��R�2*d=�Z�O��zJ�L�_#(� ��Kk(M�*Qݗ&b�I�\b�0�}�rR�sY�X�9���T)'��s�
�Uڎ�쿺rAe�N�I�(%7��+z#B���_�ts�3C�,��!�4���81	�G�0;L��f��BJzfE�%I$�� �sDJJLQ�u&~f��u>�Ïj'0}!dy������O6m��J��Ó((���t=(�q�=Q�;��U)�?z-�n��?km����y�(Q��g+MM fxsDt ������D(� ,�P��
�tC�G��v7_��㷈����B����ư@� [��I���]~�(d	O��̿������F�D��'{%�cU��s�􁾃��O��#�r�X���1��J=�)62ː`��D?��y�'�sr�<pJĲ-/V�] |�{�%���5�oO�^-A�7/�5���%h�|Խ�:3^^䢩�"���o�MN)?|оAP����]��ƤX8��M�Wvh���J���ڷ�Y��rH��~9w>c�d���{���g��ǥ��B�xLwo�	�u�;'�� '�p�W�[�3�G}a� � ����Iwl���5L ���#Y��<kZJ�8%�C_�p��f�C�c*�N*g������	{�F)o�?@�D7�F[\������6 �~�'t!�>����w�b�>gLy��#��z����e�5�jK�+����,	��'���2Mw�mz�r��V{�G�����Ccz���:j�8���~=sy�#֧4��~K��J���7�O�` �3-�޽�� ֓,N�߄�j���K�$���k�f!R����&/�M�)����3�%gA+��TS�:I�%^kIP��q�����J D??zJb�}�Z������2�T�X��qޑ��3jǗu�M��� �ׁ��M9K��R� +��Eg��e��D��NA��D�&9�狽���ƨC���*T�sSŧ�!��;�w^Sz+ B�I�c�x��/9�z��+���K����D��Z��t`�-B2'`x�2�S0��M���5����:/hK��5s�����m���
J�xOP
�v�C⼾KBG�/�*4��c��mM�#��r��M��̝ ���-*˱�8V%�˧� U��\R�q�%��u�ʒ�<Vj��|:�(og��\�ȷ~4���R�i�!����9�%�[lӲ
O`7ں�O�S꘥��~�U��]�y;<�D�T+'�LV�z�ȑP���g*�璲�0ă��5Sv�͔�j�MϷ�����aRp��I���Xt ��WO>��aJR��B��0e=��*�zُ���%o�$P��8`]���%�5`x��٬A��}�bT���k�8A�K:RL*��2_.K���aZ�B@���L!&�^q�O9e���MAd��4c��t�<�!��;>8�(hkrM�����iC)������Tm����s1���L�*)�c�&�
#���`�\��0.�$y���