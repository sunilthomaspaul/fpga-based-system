XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���"��)JwQ��B����J�s|����{��o`��H1#�!��F�a&Zu
He�K�M��e*Y���?�܀����ҭ-0��g�]��o���y��a���w6p���N,}�^�vHd��	��a�J�j���Ckh����|ӢVu��iZ7�ܹQ�3v�V_��Bm��gX�H�B,u$չV�°�mP ���r/��^.Y�Oko��ڹy�ܚ���e�m�Շ�c��\e�p�(1YI/XN��bß%�����&Q��U�߃>Ǧ�� J�5���,�P��?�ne�zns굎}��	��^8�+���p\ ��YK�E��Z?��@�h���`=�1d�Ko0nQ=���4r�|���Z��t��B�OJǾԡކ&3��Z��ɓ[���D8?�+�Jĸ�Qv�}>cj���{�j�%ؿr��d����
�kv�/��YJ� i��#�W�5$���5��qb3����طv�z�SUZR-��e���V���u��}�+}C��-\z�?��g_~�T�#�@�9@S2������<	�D�F�R:?ނ�SG��-h�N)��H�?�z�칞���e��C=�P�f�f�v�ޥ���m�
O8���S/���~�p�Ϩ�G�i����N5�ɽ?�=�'��˽ɬ%gR ���C}���l���,#JX������&�z�|�[q�u��u#����*��復��L�����F{�y0��M�0��W�md_�K��4R�k?�w-��Y�=�9���E.��PMMԂ����4xF|�XlxVHYEB    6ff5    1760�?�<h(�1Vͭ��Z�Q6)�*����Gy}ŵ��s&��u=�W�{Z���q_���<����1�k��Q][i�e��D�l�]��`/��h[��$�n:���<���B4)��+2`ب�*6��%d=8��%��y{}WAp�Y)l~k��^^�zF�XC�#�dwԁ�\��\�)��C*�������̤��"S�~��i�Kr����o92���p���Q��X��i�Z.��������|=jJjM^C���U9�&��;����ǒ���}��}���؝�j�#�ʗ��b+�j��^p/;�w�K���4�����'Ȳ�f/~��&i�g��|^\��p_l)ˁ�&�������k__�>%���S� ��-y!~�s�� ���c\Ӛ���l@{�^ð`�K6�ԗ�5��~�Å���~p;���;gWv��L������Z��C�_��N�~��d7;�j��R7�Ó�WʑY�҅�&lN��h��s0��C��H�^�1B��u��硣-.���m�\�V�ȷµM��r��>�Q=���P���xA��(�	��|z⪈^����q�)�&:����!2?C�[b����x8���V��<T\���5�n�ZF+��{\L�J�-�r�=zgF�-xs��R�Nxmy��:1
O:��,�7��H))�ǈ����V��a�����<q�n�/�f��&;@�0��:�b%������#p��+���xny�˨Z��*
��6i~4n6�&�Y��0��/%+(�����5[!�}��Y����b�����)1$�eRy+��e�0��B������^������`��>E���"{O�����<AƄ�\���Q�\�Y��W8�m>�͚dE��G��v��-7g���Er�����h|�T8#H�~�:uv�hv`�SL(��?���l�r.ޱ �t�0�400�Utw�������K#�b2��D0y�A�a��;.Ћf��7���dZ�z!g���!��y�[����_VZ��� r�4�/��B�`x��I����N���(xX3Ni���!*(�� &"�0��b��f]�݆�w&xf} �ʹ_ ���� ��\^7*D% �"iY&����[=�8r��0`�v�"�Ǚ�<�iW�p�<�Ey�gϽ�R��}+Pʰ�g\�Y���e�v�-1{�F$��d��0�
���.�|m�3�#A���?n
��*����5�|y(-}�VK��s��it�(�y���	�L..��D#�*����X�����jDT>N���'��F��l�tf28�!\�	��6�Y������&M��!x����U����+˼4v�ȝv�$����=�F���n�m�DN7�2����P� `7(p��D���<N������m��T��2#�1BҎsA��=6�l��ih�F*�����sA���.r��s��xr@�:j
�i�Sbr6����t1G ^S~����}�N��N3i �.��ϊ�~������5���-�~���k�V�E)����m�E�*	c/]�'���\8����Nw�%	�8�<ى� _w4�iP�E��yb'�	N8��(�����>�H��u Wkz�y��(�˗+���>��`H촆����(��y�����B��	�^��������CU��JI�� _؈X.iP��?��,bȮ6U�La�j^�q�/� �2�b&��ܽ��l6i.�����Q�P���7Amlӽ���0-�6�Nۿ�"���0��Z�<���tK�Y����|1:ƽ�8�����������n}�6���R�f�w?>SB���붥�ӳ�ӥrf��A}s5�U�N������Z�O������l��l�4�T���O"�ܥ��hn/L�z��xv�b2BOP�9�Q"�Y8U(�B�"��k�Z=�Ap'w���Dd ���޿Y�>Z��o�![ �1n1�ve�rb  P��Y�����Tp� �_HR����s��g�mPa�A�f4b@�f[��n���U�|�c-�i2���<��^���k�ȍi0nث���j"je�zp]�׷��vڟ��[�����Ԕ 7A��:�[~J<K������'H�^�3�m�sk��\NTJ����%l3�
K6��^4�lדZL���;��@)�b�ܸ� .6酛�H4;-t~�l-�
"�J���^���<��鿁xj��	:��6�H�Y��a���{F�� 1$���m��(:�>��fW��J�%ŉR�C��U?�cOF�_�T�a͔6�DK��tg������YG%�U6ペ�*A������.�����	p�H��h���U�R�/�8�elp})�VŇ=���˂�r%�A�WT��-��A��M�;H�< �Q{�o��z#���d;�gϺP�N�s9�E{�񭶄����MXP�O�"~��_�p�ۦXyle�~?^v���T���������Z���|����J=��Ai�ы��)�~�k�?٬<,΅�+TfK�Ϗ��E���k�6�o�t>B�39W���4����W�t'�c2�L<�i�&�Úl�O!��三��qh#�	����|� ��)��=uWFYfj60�z�yG9��fsz�ɊtbhG�����y*{zX(�W ����c*1=��}
fV�>Sk�s��I�3�kb��t�&��(T�A� ���L���&���)HN���(i�p�͹&��.��\|ʿ�,�i��ǾؑȈ�c�f:�~��nҕ�"J�F���9YO�>���i�E��O��?z���z0����f>ZN��?Yt�T��S��t�!H ������Eʣ��1�5�� �3��?倯 ��cL�)gҟm.t���2�߱+�� $1��)��\\9�
Pσ71�i﵆�'�&��)��`��e���eYJf��6w�(y��j4�g��S�2���}�&ލ��_��T��Z�ƹ�ii�yDÑ]�^UG����y�[?��:����\���w}k��ĭᝂ���7�i��zC6�#����������;�a����sQ9$�J�)%��΍�(�k�a�տI����	��y��"�l��R�%l�/Z��.8��pJ{�<8T���I�9�@0N��Q�ӒC�FP�X�yC���9[�vT=��<��<T�jJgC��Τ��g�9M��x�⹣F�͒�"�����+G$��U��y��
}t_}�m���C�z��C���=�ᘭ�]+Ig�U��.�&+,GL�����dب6- �3],c�ԇLG����Y�t�����t�v|ƪ�2wD�/��k'R�DQ�u�i;��SF��q$�A�_:T�.�$���s_������RcQ�S�;�n���)��d���ĔܴS���U�Le)"7��zJ��Q͈#g��%�C7X/�K�r�  �*B� +x�59(���̀�B�"�&��9���C����r�F���z�R�[��C?�B��q����-Z�G6���i���jD1���~�
i��PΪ�>�Rso���x�C���_g�lp�)�Ɨ�`��\�Ũ�ҝ�!M�W�,��'񿬠	�*]n�0mGNÌ�rI���	��������	)9�|��h������!��Hh#"NL�4�GC��~�@!�6��2[���s΅��	��Q�ǸhUW�6e���K�S��Ģ�H��ӥ��Q!2X튡�Y �)����*u��7s�ŭ]竈��AΠM4��;�~J��'c�/T�)+��� *���kp�{ ��z㏚�D+T����
L�۪T�=k�:�Gy���)�:+b�OQ�9���4��@5\O��|�L��U���p]����Vl͈�&��]�kM��� ݩ��x�Id��L��`���@p����[J��=�kM�Û;4�������(�����jm_T�-
�
y�S𤆗-�~g�RN>�ҩ���bu�FĶ���|J��XZJ�j-��T�;e�g�����_��}+�v5Sj�M��Y�9>Jx_�ҝ�ޱ2h'ƿ����n"�h���l����$?�O�9�WI�C�K�/���x��F��h�GH0E��"\��hV����lK��Xa#i�)������6���ԭ?e1��>�Z%�v�4~A~6��b�o�Ht��!Z�ힺikP}���MU�E���N������΁C��[(#+�K]ɒ�c�h%�����|o���|��������?�;{�[�J4wwkJd �^���AW'�'"�H��|`@vԎp���CQ�����e���b�%S|V��X�<��o�V儉�=/�Q.����V0��_&'����s���(��}�p�J	�h���/-h,@G �{t�@�9l�G!p����p��L�(�\b�4�G9�e�~�3����9$I�3xh""v%ԉ�^C��0�f)C`�#M��y ��н�XpS<�y�_�߅�'��Ͳ��^��vF�m�Q��^B�ꊸ'ok�H�I��� �<WA$�ӊ����~C�`1�����9�t�c�p��/|%���_�& �j�ٍڒ�i�MV 1�qsNQ�i�퍓�+u�t��ΧK�<U��ma�?D|�%��υj�
����I�ȸ _�9qy�����*���</ذ3�h��P��l�]�ױ���~�5R�e@������:�%�����a8]�5�E�������V{b���v�ޛ�0$�/*��	��
i���'�G����cq�:u�/B��h �;O�ֺx;KA�-
���b����V"^���Ź��2߭�`��|�`3	ڢܼo��e�X@�� ���o��8��G�|%��;��ʎ1ce��;0�$���H�+�L_�&/��W�����ѵƽ����~6:�ʎ�M�����t��;�9����x[^0d�k=�ud8wC�Sנ��$��`���J�ﵤE=���*�[���)��T<��i)���y��MNo�A�HJ�R��jԀ��0M����D�f\�/��_)������f�>T�C�	l��f�W<(�<)�uKQ�2�y`�m����kE�m�?}��^��[1����|EE��8Z鑑.,�zdD��f6��.t���H4�!MX��&2��������pH�L�FK �L�ݨ�&u>�w�����]��?��xt�F����1�[_�+�3L�wg;ߚ�DX�9d�Ym����_&l�
W|gh��w�5X���W�A8��d�)���к��9���V.��E�c��$�[�8��<��m�6S���a�4_J�M��@8�Q���f��I<f6�1"����Z�E<�F�Y�b�-��B��m,<�_𶹀j���XO{L�LՍM�b�a��2�uf���Br&7�^�f,�OT���ػ���P�;[����U(�����n���U���\�V��[p�VL�����_�}5_�PQV%�p2���&\p�p��Qn8	�hR�.��+��ϭU�:�m:�Z+sc�h�O�*3��F˭Yo��[��l�X8x@U7Z�g�Y���)�nꉆ��q~*H�<'�����&'�<���R7������s��_��y������/��+B��`
��� JYy�����&��;�����(G	H�MFyiq�u�T&���A��m_�pS@옜�b�tF20$KŚ��آ��erM{��ea�%&��z}��ڷ��QVf���6�Р����)`��ǁF����,� ���\E&�sH��G_� XrY/�*�������o�2$>X4���T����=D��;�h=��1����T����YP��%�9qz榈��c-�G׷�8�?ȵ�O|�c���<�N�H.`yr�.\,S�İ3�����Rw���#k2�
�O�M��