XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��w<���ݵ:��Qö���P:�[�7n���]G��<���'������C��˞�� ���yrZ1T�Y'��K,�v6��H�
����J(�?gS2���Zf�"l���o�pl�8��j B�_���	w�k��;b�j��cH�Bn��MQ NX`\OW�!�q6M�,�/��4�e03j�3��z�xዱ7����o� ����*��11���Hā��L���@J-�B�Gz��s'W�K����)z��*`�:얇7�X�����*��8���h
9Ò��HD��K���$\?�.,�"�>���0�VP�o[�k���QS���F�'�+��R�P[�9�_�� �7.�Eo�z�s�K��'�9�R)�_,@�7'o�*^LuDWj��n��������r����nƒ��,;�y�b��J�$����ٹv�A� ��PL�˳6@�H���K �� �����2N3K�%����N�|�A/��]5u;�w+W���"_������ƚB旎�U	�(��-X����x}]T�����L���4�'c�֓��x�S��U�B�B��/��Rw���r�kگ���c���X�m�4������ �a����H�^��.&��%�rr�s��	2!���l�yo��q�9��ć���I�nme&�b�����Q�DO(ߏ/��j P�If���:'����@�\�Pc�S�h3�{(�o����n�G���g����#%�z��Ji&0v�/���l0�\E7�cXlxVHYEB    d81f    26f0����;�����5��1�c�6��B�/�0��M� X_g���?u{/�{F���k����{�ĄGz���t���l<U*�!"O��\�AA~�G���Eg�=�]�v>�[<�������B�3�^>�+�sF~�*+A0�O=B4����~FA�r��d�h�(d���u2���)d^�� Ⱗ��ݧ<�z���̐z�/��X��:����T� Њ�����fp,ɭ5�x�����T&�0)�ճ�b�?�_��O�0ܔV�#ί�wcOQ<�;�H�����l�$�wF�ca	zj ���}V�������"��	CdX����9��	�DU�߇����R��+�iT8���!���z)1!���Oox�e����dYև�s�aj�;UL'�O_��I�ZK�� E 񟕠|J��WY�ހ XQ���Ֆr������ڵ�s����Hm����J#@D�U�	Ɠ�d�%�����m�<�(lIw?�(zM"��� 2�Z�V��7?��`����Ƽ��r�tSl9�S��f�詞R�+!��nF[X��V�-'!�qLx�b*��/T]R{�HA(��=�۽繚��2��FK7Uz�-]̀�P�R0\Dp%Τ��N2+��d��d�;��z�:�-!��X����&�1"�1�ȗ����|���$��<D��mȴ9k'	�HN�P&�����;C�`(g��'�[NCN�D͟kwt�yD1X��/5� vϖ�x���M'7'H��uB��D_���6r�;���p�I��;���R�"�h}��g�o����	Ò��&��,��sD����	b�7�^�� Ж0t��U%M�1��loy0����(J�|U�؏��Aa}��bRʀ1ϝ�'1��ѶR�P�?<��Slr^lݷo�v����v� �_Z����%j�I�R�h�2��Vj���:�¤��sv*�
�1]�NV���\
���ɕD5FXu����iaS�18(���:��x��н�p���L\��Ww����t�z~.�h���H���vb�)/LŬ`�}N
�o�� #�l�&y��'ί�c�[�W���i�� Rw��P�Jn�/S���m^2aJ`2��t�p"�I$^��HI�B .�D�A�-��
��@��Kĕ�-��D�z��+B���zK��Y���il���n�$bA�F�He����	��-�0l��zp��j/�_��^�b=����г�3mY�K{:(7���$"Q�,��s�03�ht����������}��X���p���А�]G��J��K�cc�K��-�u7:��W@���z������Lh�Ig��I����
�46��<#��RkD����AzQ���N�(:��z�c3 `�LT�|�i���U߃�
 ��(�DfjyPY��]���ؿ��6W���/��,i���77��Cbdf�q#[����ޝ�Hko��z��ٹ�6����TkЍ���R��h���s�y�&էEg���Ϲ����|�`w{�vgL��I �Fk�~��V��%�LПgW=f�Zm
h��=3d�t¤�yo�g�w~��֓�}����+�M��	5�7��QN.bHbC_	̊�07e�}����>�ot�__��bg���{��(�IL$|�(O�w�#y�����������{�w	�M�9��YE���Z9�WY�R[�����`�L��a����2�����P��WF[y���UD����*p�9��ܔ����E!悐f�]0�N]�[�Q��B��;.#D�m^�x�ע4���iۨ@N��2W�X��u��,�w�C݌x˞�0�u��}�v|�^N}�kD�f����H�,�p>�O��k/T��ሜi��XgNg�e.�� kdY/G�жs}#W�B�ގ�H=�vB�CI���?��v.{�,�GxNY�ܰgwc�w}�VWV�j��φ���&4G�֪Y5�b��Q�:���i��ڝ%^}�����W�#\���Wrv�r-��b���px�Kń/X�)j�
V�ɯp4�ck��^��RV���?|�F���@ei~uZ�g{o�X�=�w  f'�yr�rO]4���7��6�)J��V�P�0��pԞ?���A&��sE�U*�� L�.|�e���w�]�^RF&��z}�n�c6bپ{67Ț_��#h�$�=��G�^�f��%�N��o����="63o��n���ƂT�k��}qU��y��G��Ywu�ٺ.��sI��n��`���8��^�W�}�'P0K����U\�<M�͖ZE�d���ns�Z�aO)xs�2�C1p���G�VْQ*��K�+�k&�>�w�e���gD�l�z�]~m� j�C�ӲƩ0���|<~�O/hz���}�֜d�?�2)�^��5�X�����%�d(S�a���u��/�ȴ�+>���3Q��C�j�ܫnN�F����2�z�.?:Z��_9�/ׂ_8 ����FOwblx�lB�|����:C�u�(�E���ձo8�*��p� .?!�D��sP5z��թ��H^�r\��w�}���7HNi$�_�f&��V.p�@Oâ�q�DRCjy_2� ������g�?"�W_�Ff����Hm�1W��$��8��W�~
��Y?̹�}/4$��ɸz~�CS�n����&�>Ne揔1�T�w��j��E�p޳�R��F<���덺��7�6c�w*F���,�Z�����wWa��d�٬�I)`Bī�����=Z��rӈ �k�Ll\�v��$+y\غi����P5r��J߳�(�����{z�[9K�S��&��Tt"�w�k��3;��x��D�[�[7�Ϩ'tJ.a��`����Çࢊ6WWO@��Rt��]tҪ�&��[�њ<�������n�.*0�z��)������S��"S���[�)x'n�_w40W�5K>Ɛ1��l��3\3pdng\H��-4V֮��I},�g�A�T���_~�pP��0���'����z��	������8��N�YP��	i\��8鴤�$t+M�gR��IHG�Ks���� .��C3Od�p��[���{��~'�b/aL�e V�%M�Vb7�����4���,�0��������! �/9��݇��M ��A��lei���G64��K��u_��n��6���s�ȳ 6��Ɔ��Bt�Gu`�+?�_����e���V��8�u��/Ѵ�*Q�^����^"
Qp������k�5����Cz��~~�5�x�aW�̗�h)۷|��_�Mn��CH]�g��_�]H�q;||��%`��ѹ�	y����ʩ�(�|T�:���щ;ۄ������+i�a�S(g'�L52�5��X��2�@����O�i��U�]�~g&O��#=@�(N��MȞ駉Y]C ��m'���ɗ���f\5����od������}�`�V�7qh�m%Ǘ�a���o���
�r9��B	��ɶ��v[~;pnG�}}c0rڳ�n��6^6�A�u����9N�A�)>Ǆ���(��u��2�!�1���z��XL�����S�+�͹���t�W�I�l����H�E������4�tj4Je*��sHNO?=Iy5ɡF�bv���[B�:�r3OHL6r�.����0X�~(���﯈�	R�D��Ȱ�Kw@��K�$�
�|U�'!u^,KJf�R�i���X�{���ˎ�7T��:E��΁5���m�~��+X����|�7��r]+��<�Ih��[X�bY��kDj5Zj<{���b��̰�n��,YyC��X?����h�)��.H�U:_+��fx�PYtS��_3z��8I�X�3d����_�~�Lmф�-���@NNm�	b��0+y���u��xB/�i�%Z"f�)Y���|^Pě]�
A���e#��e�Z�W�����������-�"��%�������)���T�������	���࿁��No��R�w�>�P`�Ct������������/)���Y��2;�e�Y���#�@�XkA����2j�Na��h��Q5f��x��c[ڐ~�Nڮ���!��%��b�W.�7�����|����G�@�_)�I&�ʱg��'�?�3����������y���o���'-��*�T��N�E"Ii��O��2�f�]�|��f�\.h��h�4�h.?Nb�{�#�򎎊Jz�J-���,go�ܠFou��M�����v��plㅜ���N���_��~�e����}�ܥb�$��� �!�/j����l���"7i�/�Q�ݶ�W-�]
��KzN4�5��P��U�Hc~ �a�]���{+aw�-�(���������B�E����"?�����q��i�N�_u_ n+ARb������ ܾ�f�a�o�͠D�d��j.�At�!!N˂�"��,��'5C{9s��it�I{����A�z���Z�2u㰦�1q�$�F�Y�4e�FIR�p���t=3�.rQX�J�T�YR��Kݞ��حa��ab��f�h�mP��_��&��!Mk,ө�+�Y�[�j��c/�؂y]�d �k���`��D1��b޹t��"U��@��n��pZ�f�<Z�`����G���Al�����T>]B����KP�O�'���o�t$� TI����9����ם�(]��	��=HGJ4�A=1�ѮO������q ��Rr!��������PGF���ڳ�ʼ���*�3�w�]�x:�����L���(5�P"��gɟ�8�yG�:P��~g����o���w��P��w0��y�Ë����Y���e5��!��� �S1u:����c*=o����l������I
�D�(9���L�H�aG��7U����C��Ȫ��'���a����;Lqu^)�E7�i-�]P:��#.z쿌"�鸉,�S]I� [K�HBws�b�ŋ;	zK�	?Yo43U�����
Z$���!� r���ԯX��¡�90k������hc�>�<;�
$��Þրt�3�P|�C��!��Va/k�m���)�M�覫��nc_"��bR^# ���jv�2Ƌ��?TS�Oג �/�j�#
����k�-�F��*)�&`��d�s95��ƈxՅ��q�&Y�H�]<)�<o����ɯ��e��kK�<�Q�����=C!�:5r�ck9ʏ�,ɰ^@�2{F��y�X>!-w��>��ܑ���x5ƞk	*u��Y�SF7�-,�_��5J���.2��@�s��Q�o���p�O5[N�*F�%4A%Fg����X��%����{i�2p�߼s��i!��Ѻ� ��U�+��V�gK�K�����'�k/)+����iFP@���%a�I�N�D�W%�~��^E���vݵ)N�F[�'�{r�yP�o�O�IQ��K�hL��5h���Sorl��*�.�F<:qO��a�(դ�+�|ƈ�Y3�����{�2S�9�`nHg�3������&�		���څ''�F@���3BV˪gHg�+a�(��|�'D���u+>fx�sJ����S}�3��E�I��h��V��t�;�x׈�I2o�����k�,�K(�O�)q�@L�z���Q����x���-;��߄H������l�y�E�q���r]��`�!��.�{;c�I�3>����8nI��rO��H�B���d;'"��O��*��������m�vcMZ�].Q����:^�!㡽���f|)8���y��g�������u��^V6�7���ҬZׅCR��頝�ߌtA�%cmP<�~�W���l��e�:�
m��̃��Ly+�Y���wo�zX${مǫ�����T�v"=�#���o���޷�4�4��7�uS�&!
�8EKp�2CF�>�guۿ��{-�-�J�w���۞���T�1��ӻs�(��Pլ��J�oM� C5_�Y �ݮ�>_I��#nm��(U4�b�*�$���o��}�t���t�-w��S�(D r����@�����|:�����'�&���� ���O>�D���')�����8ŷԮT:���׏N��Oʬ[:"���pB��t���/����X�v�:��a(�ɥ�"=`#�%y��4s�CvJ$۱ef__k~������X�.�,V��7��/���;��a�0��`�����RG�-7�?���#$�?6rW#��"�H5YN��3%�&�ů	��;k�As��^�(x�n2��}F��[m��D�Nt+ =3x�'Τ�	8���l'b���d�j ��o�'��۳v�E+�� Uߵ�!���\ !\I�7�!��I�2�./a�����[]pF7l�[��ӫSw� �ޫ..��O9��A�J���`��}�}.�Z�2�d�����Rb��o���瘹��ͳ9�NZ)Gx+��Jt=F,��.O�|�īM~l��.,���9���Y�sn�7%����s����nV�9JC�&U�[�X�\Rډ�\�O�#���A��3R�Zt.Ū��P'����`��j����3	X�s�|��#����C#����;����za}B2��0IXi6zK�����if��s�
�� I�#��e5��N,����(4�g��$��|N��`�z+���i�Ѐl(ny�%~���;�^�iIh�������-��8�]3*O ��`�뻑�N��*��)�&��&��'�kcQ�۬���p#�rD�Z�^[�`I�M�Q�}(I�/@i��cیR���IN�ݳԧ]�x��?;�1�o��{�=�9�"���6��v����:�t��?�0|�3�w��pG�����Q���X@�^K"���L��,��mssǦsx�H-�D	e=����H���:���f�M84���ּ����U,����?uR�������"',�w��6_O�&I�z�a��c������֐f��qOĶ���=�0m�cH.鳮K�S�L�����F���(յ�,��i��G��{|�f`�(s�6�qR�^F��*��}9�1h�����iICC#��ʨ�v�3?�/�<�w-�łC6���C�m[�WlΜ�EH�ߙ!°�߀��~���ۀ����Tv��s�\������T�1I5C�yǎ6�:�>��:���U�[�Nf�y�Ta�͖�r������i�x��lG^F�5��[؝D�i3�`�Q[򋈠�@�l����Q��?�-R�Q�Ֆ���cV�����~z'�u���w�<Y��>�~��We$���Ra���X���-��:���>�߶�[�sZ���]��VW����E!��96rC3�H��;O`JL��g��e=E:&��FyiH�|�m���W:x�Ǹ$�ZL���ҲT��p���E�@ذK$`�'"_�&��tG�o���DA-:ڂ19w�r�P�}�dK�A��{4�s�mV��d���%���Áϰm!�������j���&��(A�k��,�*� xg������k��\4�Ft�6�5����_X���*X���FP�D�u�P���W�d|H���*�w�7a�h��`���@�L���s"���L����� ���"�<�ô�����zm�E��WA�l�֔[�T?���\���w�h��y0�����t��r�|�ة�<��۲�jʸsB�z8�3�H��i�����I��G���/HYfL���]���e-U��Q}�H�<�Y�JI��DI�^��rd��|`U���2�(��,�m�=�\~݂���;ڬ�[Z�^Psj{h6!��߈������8�g߾~����w� �R�w9/���VE��^쐬~�+�X��Q�R�G�
�S�싉�+��)�g�܆�]x�/����y)yF�2N�@��!��S��
��	4nZ��ńL\J�o��E�� �J��.E�Eqm��a�.������Y�Q8E��,mk��7��
� ?�X3Ϋ�a|z�.qsW<�S���ގ-|����=c��������B�J�z���!��u��h��)��i�M���2��g���#�̓���]�S�/��/�w��5P�3c�[��0G���B�}�4�'�|V�j:��[|�~�EtVQ�����w��E#�v��֤��@�!���k5���<X���J�86zB�������J�M	�C�*̴��H��Jp3	`����ZL�iwh�S><H�����r[�-9�T�[ _�lܻ�����Jcs	O����T�[����+dcv����D�R@2�̈́Ein��@\�V{A}����V�7|/n�Z�4�͜$l���/�Nu�{��xH��H����\��S�X-u���;e�U��<9��+�+xI������ \gj����u&�dtc8��;&UC?��l���c鋾�4#�t�����T�M�6�������T5���ό���z�-#� �c�o�f�}�4J!�A������$�K_3a'{^��P�rY��� ����<g{��&Rp�k*T���8r��'�$��(������ِ�-��0S|����1,M�g��1(�������$���*4�M
��J���Ŵ�AG�WU��vA�h�j��;����͖goǻA#��@�f��7"�ʁq�ٙ����2��|'v,�BU	�;<�մ����^��|�&f)��/�<&�2��]���3ЭS��giƅzv�7�UȔ(���c-\j���Ά��pqN(���wkn�O"�8��d?p-����=��
��d�����xt��cJ��E���y�[Ǒ��=>�R�O
��n�A�ǕŇ*�?�	�L���/��X�������ϑ4�k؈Ǌ����d�é��a^Y�/e���q�c�چ �_�[��	��ɜ���5MM�h�eX��]x����B��oX&����V��~�U;-���0@�E�_�@�AFE��c�����$U��������|):5m��^�I�j��^�5Q.�A
G
t�r�{"�^���n6��E�K��Ǽ2� s��rh�������d�*ZN��&���(�N�����D��y3w�JE�U�Eg̜M��gd��g�U�1Mfrr���!�u�U��d��KB��KҧY������.�3�-|x;�6�$�Ӵ�
�q��W�	l|Q��/4����d�"Y�NJ�
�J1ܵ���^v��0P����̚���bz�sд�L��?"v��ǀ7hɕ�����w��n�T��"
r��y2A���ަ��mLZ��O��  �nuJ����gݼ�	"ɏ4���{���dXp��H�Z�9 �|׉�/���[�;t�>)F͢�h�U)�]�Ӯ>e�Ome���	5��|Ń�uK��}|C��`d�rXB�d�B�Lן��$����@/@D��a3��N�
��p��s��ۍ��}��k6Cd��tT�����͝_~�E��0�HE��iռ|�s/����y�&�V"m*R�5:��BT�_�S�������z��\�%�����}.��m!r?*ߧ�M���F�P�j�
�:��TKC�x�zt/j��1��,]���֨�C��o�VA�Ad'8�h;-�پ3ԓE�������fEV��
$S�ب���Լ|-��Q���$�w��`k���R(|��Ok�[��Vxۘ���7eiP����
����bi��Y�U�@��﵃��k�R>F�����mw�����Q�N�VBC�+�.+Zx�HH�@�V��)kg�?`�$�f��F�T�yFj�ku���	�-��l�	��TX����yUMk8��