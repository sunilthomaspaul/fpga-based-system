XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����O�/���B��*��w��WX�P�C����!�Bǅ��b�fZuP��w	� �ܓc�����T��)M�v��'tb@[܏O+UKCg`�X~�8�+����]�]	�͙g��
��ȍY}�u�4/]*+�h4F$�s=��W��Re��ح���HMà�󈎝�y���^��`��v$ҋ֋À���0}6z�y��O��%7|�����Tl�5`������I�w�<�]V�lg���>�g� �n�?!��Ub�E�b+g:����X�K��o�Mx�P���1�{v�H�l|=� )��i��?C�S�p�ҫ��͋3$�Ȍ�>&�� �;0�ן�r��9���k�@ܺ��A�q���S͞煍��L�8³�Z����7��vT��ׯpY�н�.�h��V��52��/ҟ��b�<-h]+!�	����>�����gqu��� ��<F�Ƞ�ʾ}��M�6΀Ť�b
��-�s2�U5¾��B`Sk`��0�Bb҉�,��~ x�%H��Tg�ҩ�~ ���t��w�-=W��~��|����^>��2�W�C	��j�1�P��욷a	(^y��8��I��u�hQ���RZk_!$�FlI�T����c���#�&�>'$
e�*7b
��H�Ǝ�m�dX��\�K���G������%��ø�q@�+�B(�_���}�*�5���� ߾�n��v��g�9��o ������K�����E¸F��,�@F���KXlxVHYEB    523b    1130�����O��^��X�Xp
q���[BO����G�y�])�����h�����a��!m���,=Z�m�F�߳ۖ̄��:�� �7�SgGH�_�ί\h�yv���d���^�AqL�K\{�X�ֵ$ٟҳ�@9p^s���M�Y�O��uCĴ�p3�u����r�O2�)c����NŖO�:��c37\�<�(��YVOuco|	XH����!Ä���v.����vg,��1c���{�sOі�܈�!]��g�S���v�߫�`T�w�R�W�%��)ۥg[�`P,�ɚE����{+�����K�� �xd�H�UW��kPF���$�暵-o;�H�K��蘖�b�~���m�	�o�0N��͉�����\el-��'� A�1L{�d2#�J}�+�D����^x�� v�G9�������sQa�a4�����E��4�Ғ��؋h�`༲E�p�s���B4�8՛mȖڬz8'"^�t�6h,A"�����@T���\�������  YV����z fF�~m5���;�w"r�Q�-�5~�I�iPG�h��B��(8PV`�T޶��j:�?�^�o�8Z�����Ԝ�~S�GI�Ujd�P�����|nt��
���+P�Ë���2�K����u��t�G,0e�5�%�E�Z���? ՙ|e���[�9%�4���n��U}�4��uWۛ�*���Ӧ,�8�{B��ܸv�K_[p}�!;�@�@��"�E�|)��;@�%y$y�[#��iIv�3n��7�mk@TA�|�X/-R'k{�3�}��I��ҫ�9;��J� ����ƌ�k�Y|�=!t�B���_������nx�Ɉ�s��-�n�]	z�2�>��D���O9+�2��G��I%Gh*��w���,h�+`�/��\�U�����V&�ӳĔZz�|�2,�Lb�}�fp�{.��s=I&
���],��(ִ�L�щ<�ƴo�}Jse�rls��ǔ��t�m������o�9�+�)w�����Z��J[��q|�]�{�U�5���c�J�)}���L�I|�R�u%�jy�X�uyp�MAL�,p,v�?sݒ9�If'���ͥ/I�%�9�П�E�wMK�VI�?`#�}�x� 8�G�\��s3�EQ�a��'4����H��6��Pu�|��S[I�R��z�<�M|md#g,�������"�� EC E#�ρi��Z-�Y�͈�V -׃�{鵹�G5����.u��4<��� �VZ�5�5�Z�p,фTL���	Z��Qס>Sk�G����a�i"(̛����o+�(p��[U������M!LN��x�
���9P�Fg`���A�-���wl8?��Z A�z:澯��Q�39yŎ�Ȉ���;���L%�����P����ή��r����몰��`/���Pc建����dDϟԘ�Wy��@|LCg���M�
�|C�-�9��H�1&
�I�G�^�S-��A0��xQ�rŅ��P�i��e���K��a���0�.Y�[�p�%G���d.�䢛'"�^ǝ>TFn��aK��S�� ���!]e���*��Lh��jWz
� z�T�X����t�h���^�c�A�&�1��:X
�����^��p�]�ͱ*���g1:�؋�i��J]�j��s���7,u��N���Ħn�Ɛ%ʏvԱXY&4b��`'�W=j@�Y� �	'q��,1S���G�[XR-lW��o�S3���Tx�.(�}���y̌��#�\�,�7*�D�ٹ3`n���)��|���x�G��$7y���ӻf'���t1�8�ԓ`�o��0�<��(8���5���}�?{L�#�S�(�j�g�]�6���S�,}A#B������G$�^�Z�n�q���/&C-L-K8BE��	�\�#��
��"�8Ԋ��T�q_{)���%$�T�_�ǥ)a�k��yt��_��=���I��D�����,)�s����	$�F���r;!�-�"Mŭl�Mh@ �%2�<ސ��֎�9GWg�Q�~>�q
��?�Pr��ڜ�${���Ă�%x���3� j�	�C��UN�6��ퟬ���W �@o3�G�����2���A��Hӑ�s۾�b.V"�Q!BR�3
�4����D�XY�Z(S�[2��L�Ay�7ky�V�~�x���:�aSz_�ݓ��o��Z����2&����U�Άq���lL�̗�~Q�L5��OB{wM�6
��D��U"IQ���$�T���s�h�C�,�}��3�a�p�A�����s�4 p�Z�>������� �,A�9���\�"�F[��M\(�zQ�H*�e���d�ݸz8� f-/��#Y�'��J�-t�����XA'"23:r+��8'~�Qm�+�]�1%Qe/�J�� �m���X9[�o��+��ge�=�c���>.Y!vi����ːC�t���� �2��m��ͮ��#���<�)f�wN��ȇ���7=��Z1�@=+�IwD��:�x�3�P�����a��Ń����Ϩ���3/Gڸ1�,[N\�b���\�.�.�SCw�ʘi�B2>INk�}귫L*���4�9��L�:(j��'�ܣ��{IJ$�"�P�$j>,�8���e�	��$x��j���AC÷-}ŧU�NC{p@S��f��Z�GdG��v�Iڬ�L2L��q�H�is�N�����V1�ub��<��2��$Y����B���/��ֵ�W_�]�چȏ>q�Y�Sw�1×�%��R�Mߨ/r��cEr"��R��韆������eJM��d������w�@:�7����U�����kZ`}�	��NM��SA�����}��w����1q�?�(Vr�@�Mh(�����I+.X�v��嗚�؅d�����o>k��3
����=g�Z�ǚ����R�5�2��	�Tg� ڌ�_ ��J'`E�K*%�,FH���T�N�I��n�u�2�|b�5}��Y�����K�hG�s���՚��☴�+:��jt�%�}P/cz����g{Q+�+̂퐞]e��(������D��j������_i	�}�pl~3�go��Z��!�o��1�F�� �\��޷�09�%Df�v�=j1;�*�+��KWǕ=z���ށ��1�$���`b�2�ߧ���OߋtTNi���3t+��
�
�0+D���&|U�k���b��'�zf��.�5Y������A!I�p4����D�ݯ�X�a�#�:��� �^��PJ1k���ty��\�aӥ+�,�Gn:7�@�l���"]�����@�Z۴��	��*-�% O3_�-sJm�2�b
-��V���T`#0����_F$���x%����K'���Ml}Я�kq�ˑ��
v�8%��A4f�̩~�~׽�;�*_}:����yqW�|��h�Em��k��f�B`q�P�L�i�Z�R*��:Ra�� V�& ���Ns�sIm���7Tm��L��
䂆Ϟ�V��a&7V"����r���}_�hޢ�
&3-l�p[�>Ш`�DD�s�����xn���)`�Ou-0�F]���g��z�䟧�5��
k	�bT���a�pW&��K �H�w�#z	��=�ǉ��O��n}�j"�(�	���/�䇁g���qV2E�Li\���4j�H,m'wu3"�,3��ӑ�9+���%��i�h��ߚ�!̎ǣ�����9*+���X�ꕚ��@3! ���̢I�R}0��%��<^�$�F��Ϋ9�'w�%��`����Yk�5��q��h?x"E�p�ﺭ_	�P�+�#*+��H�*�����ZԈ%�e�in�N�;2/�]�Tf���m1�, 3�J�>���T� �2.��#q0`Ik;|����_3�6���>�Z'�雪w"��#Wjt�y���9 �����5*�
�(#+|���P�u�{��B;��2����������m�ᇊz½�w��T�/Hب�WY����fl�� ��Ӑ���n���X+Y��GL�� ��9� 	Zx	$)��{�H�A��';����4#�+P�ff2�6'���R�7X�TQŧ��'��=��Bh����O���AW;�Jdr�D\7�tp�F��nϛ�N�!Ul0�/�,�ȿ�͍�2�*c�$�����������&��&�尭�XQO~w+��_�d_���������¦�������;�AU��zE��Ğ�#����}q��9_����cr��^ʌ\���㕿���oS�� R�r�kk<���g9�AM6��կ\��\F*��Y��Y>ѥ���=ºL}���P��#U%�N