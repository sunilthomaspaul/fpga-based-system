XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd������<�	�Y���w��n������XUJ����#7g�� ������M�'�ٺh1<!cJl��-_��,=�|���d��;De  ��z�/�k�&�y8z���.�{�K�j(-��2A�!w�����(7���U`�j8�*����Q���eǄk�\ᘲ�Q�<��y[�f�=��@0�&0��p��p�'��F�P\4O6 �����2G ���1�e�yDW�ƨ��N"A��w�he0��jc����f0��/;J 2N�#�w��j�RC�"𽚚Y����o2��%�o���e��l�h�C�ax���4�������_�Wr�s֝��
�xz��72ͼS9�1��m�����$)��Et�}`E],o��{7t�@���:q��FV̇�r�zMjo�!����pOP�%[
I�e�e������¶Y�_������^��6�c��(�.�)?15@0�ϫe�ЅHq�R�&������h��rJF�;��6�)e���񽅡�	8冀�����	ht#�K(�e������ϯ�mfaTP_zЅqg!�SjV�*��z�TC�E��������v�os���+������o�P����Ҕ+�ubI*� ׼��!��+ZZ�yC���+�SE�)��U��x$���ea�$���Q���ۂ�.� e��i�ؾCJ�ɾq|�8㳠�QAL���Ye�{�ߣ{��o����$!!�je��5�Ÿ�̳�čf�E�w� �5�O���XlxVHYEB    9653    1860��1}��k�´��L-�"f���[X��os�X(ɠ45��/p,�D���=1.Ho`:�G�7�Q�}���$RKvo�`k��;c�R����5��)&���a�_�E5��n<�^*R�h"��J'w���6)��<R��G��0]-%�����`����U��,�MZMZ7����O���6���(����=Xr)�(b ��%�4��k\�
p@�)I�9C�ݴaCj2+��k�:̾�;��kzI�p�XO?9���<���aI��RK�Q��
 K^�!����6ф��ЧG�U�T+�	X��'ݦ�^r���*��6�C���w�?Pmm�E��J���Տ�`���%�81��i.�i(?P�/�.�1T��Xʜ0��Q����J��%�Y��Ć�9wי��'��$�)uď��J=ؗx3&}������Y�Ϯ��fo���%]��A�_5�~ ��?/MMVV����HO�\��Yq��E���;�h<	5-rG:��!�;s�m�آ�}F{0��ܿ���J�z~�C�@N�"����C
�%R���\���G�%wM�q-��v{N�T������J �.<L�+"J��۳�SG3�ƓֈD���>����OPw�$���^Հ^u*KFr�{=I�G%@&x�
�j�`�`k��Č.k_�}��$�<�l�(&7�R�*3�Y�#��&�֭H��2��vտ � j �)\�*gὍ٘�:!����*d�b7?n�kwbӭ�X&��������S�z5}8����~b��p)=�����ۛ�f3m._���?�i��������˞�q@9<'��uK�<��v&�0����`>6�B�8Ɠ�Ei4m�^����/���:�4��b�8H�WS�ye �\OE���Bګ.<���\JW��Ãv�;'�! ������֗,����+��.f�m翸�v>�ݵ��"16�äg�����O�����-(�p' �Bo|q${A����y@���
�t�05;^�nY���W�Ն㺅RN?#��Y�yi&f^t)E�G6w���La*z<POѰa�ζ��{I���?�g1<T���B�Pg`��-t���n�dz�bJ�X�X��H,A�<}9�Q��
w�Fm/DH�_X���䊳4h8S���rp��+�=��ħC3꘻=m#���_Y�z?��@^n��)N�^LU���RS�i>���0�Ƞ�䋵���h�4G�%9��1��_���E �"B{�#0L�-ֿK5�p_F�{�%�|����KxB"��Pކ�������OE�b�zf8�Y������J�k���2��	iH��WʳA�*i ?>�����$V
ȩ��X���Ey��t�5X�=ڜ�%��CYɖD)t�к� *]��]�� 8��$ސ��Ȇ��%������O
k�i�iC�Ê> ��1�\� /��ؙ��ORzL��($uw�ki�p�q�M0�����Е�o��tu����#���m��=�^��& �Rs�3��6�卅 B��W�U�DN���lɀں�������UF���!��.b��hDS��a�9�reV��M���ғp�M�c}t�iF!�,P0�S�F��ہT�O;�֔�lKw^j�ٞg��Cfr���AC����<�|�o��p4�/����$Qh*�Nb����$q��f�&����y�)���`�e��2�5��y[!a��R5�,	`��t}*16L)���2�kIv���*�����Ie
���>��j����/S5A7F��.hF�����ܰ �*��r�
q��`����Aj��wݷC�v�KK����Hr�U{и�dg#v����9���ȋc���$!��ǰ]��p�����.��=�Z}����\��� �q(���X0=�NLN(���8
�oX-���q�ߩ3�#櫔��=s�+-S[��!��I��Gɪ��a�=.��-���6i
SL��_���ϩ�s�^*#��N��fcͪb� 돃MkSi�k�qT�7�.m�¯�a ��B�$O��a1��@Ti��&�U`{3�.
�E��P�,�;��Z��A��|�b�i���m|=&*(��6(�!$.&e���Wc�l}	o=7e�7����6
��Sv�Qܘp�4\׷�,,8��F���qu�ɠ��9"���&�+B�γ2/s(�#'3��m��O��)��e����l�� ��B�W�(2tT%/�~,�c�󮨨�<By�j���uE*���nG��}��N���.~�&QV��߲�%�bAT�3Ǧ"h�#HW�9�r .�m��-[��7}q:M�d�2�f��Cҹ��,�J�̂���~ِ$ڦ${�o�10><�||{Sp�~<o7Q^��z�;����hija$n7����ˤk���%|&0/���z�p������N
�Mv `��tfL�ԭ�
[X|5�~���@�����ls���߆��>�EA��}��h��k�b�	m��z맩��q�x�EPD�0f�����Ϸ/s�;d����l`Ȧ�Q
AC�mǱ.����:� �T7��^F{]w��U?M���JT�1�}�9�Β	3�AY�Ξ��S�oD�p�3 "�v?HY4@X�М`�m�P�j&ҿ�%�����9�)��>	g���9��
��}|������PC&�C��ĻH��k�<qc�	{O�����*�Pu4 �����u�4h`W��0�T��7��:��������OR_�_�~W&HLK��c���R�KM�ju�u��dw�V3$���^��L��������+�Qأ�C���p^�?�U��+�%P?�Tɚ`mu��p��]T��;���!Ѿzh2�k���T�>HJ���1����u�Asnz��KQ�D��X�!r2�g�;�`��%��y�����i���-�0� 3"�b����~⑭C{йD'v��.>bU&W#��@��o`����vPY9|w2<�����Mv��eL�&1��o��OW�d��`��+�6���k�Ԕ�����N��ȿ	__�	9(n:���Q}I����p?3#��ι���>h���y����H�AU]�D��U�fC�\�)�CC�IP�豺{�`�
����Nx���d[L���Uo��%�^#�ٵS��y���t0=�MPc�����CSPh,�{ܦ*WY�4��$�p�m�B�3'�*�k"v����0��e����N��KXb��,}oh�U��~�W[vq=d�R_�\{_����}�lY�eV�VT���X/e�l\S����g��������o). �)��������yVP�A4�����K�Y��E8��@�@>���Z� b�1qs�t��~zf+-���E�Տ��cStSu9A����mZʕ,i$�R��C���	s�i�+���\�D�FT�<���q�,��o�l�Yi_���ꅭ�l��r�z6�dm�h�K</�� ���X��v$�]دaܥ���X�9�{я1���Q2}�!�.�a��n�m���84@�����P��&d"�p@�(���<�A��@��} �C*y�/p-��Ca85 {�<O3�����o8T�D��Iˤ��aY��B�r���0š����������o'�/<�B��zk�/�>FS��Y��8)�=fr�9����z�>�mc����Bn�����]6������G5n.B �:�}�š�m��^��+��D_�f덣��p������E�f�o\*��S���%Ў�����D<�᩿<fZ{�x���n^<+��̅����s�BB�j��h@�E*�aꏻԬ��K/�rZ|��J�[��M�ʌ��0���A��i�P�@9�ǅh��}9Kj]��k�����y;����C�У?�u��Y@��ޅź썣<3��
����ꮻ�L~މy�fƲ��+��;�Q�I� 	�x���!�h�PKIp3� @������߉�`ĒO1��]40	(�Sp�e��A����H:�e�����el>��7�g�Mr�г��H]�Q}��C`�ېH�y�)��xSi
�q�8��r�\���^�g򅐢���rg�?�w���/�n�7���̵�8:@`�6��p��0,,�'�]��[*T���i�� ���>�!�٤���؈��X�xw���xN"����.�L�E@��}��N2EiE1)�_<ω״x�b�4�������׿E�R�C*U8�D|_����2��lJ&iT�:g��e���7�X����x@+T������8E��	�C�̉*��yC��9��V���y�K����!���x�ߵ�W�	f��v���rx��}������ cBȆ`�9cޜc���/7F�*4�!+�ZԿ�4�� B��5q�,0x�\Z� �8������5v�$
chd_I��b�ô��ܗ��}ڜF�6V��b�M�z������r�q���y��i�G�6�$�tlW�Ã-#~����9�~`��	����m�
���^u>=�d�c˽U���\��j��Ѐ�OA��j����}���I_�����$g=�K�Y�y��5�>}��<ez���_�")���m��"��r4	K]!���1w`�K6�YWJ���������8�eD�HN���
��r�!!s]+i��?�����b�%�X~�K�XjX�y�p܎����rc�.�wB~�1��̇�w8�e-�B�aJҮ������I�t��W��t)c%G�J/�Ňx����t}�H�=� �gֿ���j�zv�'�k���6�����8���ܭԉ�`K�G�Ѹ��Ǫ�}f(�Ax�$ 7�k�Z��1��T����Cȥ�)����t,���(��N�d��wO!�ԩ�cK�IӚ�2·Bf�5�s�?�P^�X$l�h�0w�v��c�;l*,�-FDv��;1�8�`PfR	��(�d2�TE^���ۛ��ä���g�6���"w�>,~W/����%����(�|��ζNC�%�͕��_08����4W�3�p"����'҈��w0�M�iP��\�;$���ÀA�Pb�ߒ���װ
;�����!�D���:K{P�MOC�D53ǈ
���.�$����O�R��&�x%�j�� \�	�7[�}Ƣ�A�w</*�̀)�B���Wy����+�-�I�)Z���	���TE�2k��e�5��ў�`�I����,8�h�6I�50��SR%�^���bT2.8ѯV�����/K{��y�ݩUZ�yG���RKtX����u�@`�s_��*@����!�|����Q��?�Y#_�nY�#77,��
^�F�)�Q�7��V��:�^e�i�l�V��RvhJ���9�Q�X?������cش�����jo�	�,���1(;�_�5,���a@з�����.h=@���#�P�\9;���
nn�} P78+��6�pblU!&\�Gnޛi�OX�Q�߁'E��.�v}�=�����*��m먮# �en���y�B���|+���Ʌù�e�ַq������r��K�l���a,ՃF�%�R�商�um����O��Pz�D�NpR���ռ�����i���k���F���NPI>��f�ۦe�=���_g{
�Y�B�����y�/��Xݼd]�)#:�����jG�f�&P��O��ɮ:z�C���{��+ݧ�i�lђ�-�_{.�)i
�X�L���V�3��o�q�If�2{rc.�N�n(��gߊ
#tt#�B��hk�g��S������Ħ0�o7b�Z��Do�K_��.�l��~�	�&;F�3�\��C�~�r�\�գF����(o���hp���,�`9�5ӣ ���s�w�n+� jYg��O_��%	�se����Ȍ!B�@
�@�:
�L:a����U�Žֆ�4��x���81������j���3��h��?> ���`G0��!�C�*��&�g���" �S �N�s�g^1�jN��,�G�8��4�-����f3�@:ֆ���΃>7�ߓ�X��q� $�4����ف%jƙP��l��uc��
��.?����N�e�I�Zm5�(I��fS�8|���c��:����2pgJ�=�?>����lɺ�`w$N2�F�'�+��L�~�_��Mr�3��8�[T�CP,,X