XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���C�	���/���$(���lkW���w��z����ƺ�*T�&c���y��Tw1x?I�����=:O 8��y��R'r���ⳋ��lt?�� ��36�8�����vs�҃� �Zy��yuYڝ�����:K]~��59D?���V�Ai�R�5��t���Q���Q��"V��Sr�щ��|�&B(�k��.a9�&$�5M�⅍�Ro!���5����p��S8�oB��Ά㠈��m4��30Ƥ�����[�k�!�SW$�4�	q�2ր)�� W/�F�6X�u�9�3�(XOD�:b0�'�{�(��/�uZ�:�X�k��X�h����%�<��F��.��{.��<��\Z{��	����ː�",��2��po8u�c�⋦�1y�^p$�%�/�OH�w�[����Z�\�)S��CY^�̳����I�8D�����|{]��\�ꌈ�����%>��J���A�𻗮�����q{��D8m�VOޔ�v=#ђ�����)�L���%�x��q����;'���9�6N
��[��>��[�=�'Q�h�f���M
$=Ų���
��4�f�5F�;1�oL# ����5���3�.k��������K������ܮ�w��_����"5~�>׸���=(�9J,��$T�Y-?��K\�캮�|�����7 7ɾ*>!,˹��r ��$@e8T�S��.��/dB���d�c�J��w�U�HZ�lT���.Ƕ~|(���;�7���E�W,�k��1(XlxVHYEB    2442     ab0R�^t)G�u�<@>,��������ù&0ҰP�zaVy�l�6��C��&T��k�O��{A� cb��I�	Vށ����oMy������w�)iӽ������WϺ���k�����i��L��L�/J���Oh� u��J)�w�����d��Éc]`��p@Kʺ�g�T]&��<NIj�@�[�)�,k
a�?� S��8�M6�To@�M��-h���*�8�����Ɗ�9d��Y^���6T<�����% i�����h�LXm��D�W�tZЩFOUh��N��P-��D�T�0�u0QZ�w��Ry�oAA�w��W;}$�� %��6k� j�Ef�M�Y�����
9c�_R=���w���r�W`N�]m	͍�6��{�$�J
4]6Δz$���I{wƲ�m`'�2��Zߘ��٨��z�7��}W�>�q�J(7��Nڒb��YY��?Xہ57��l�8=%����F?r����9�B_M����@�%D#����ܬ���^-��Bk]����acOѕUӁWa���p�Q��<��y�)���_�7w&<�"b�����T��/5��� %%	c�{�@X��a��J����0h�	�C���A�i�(��T��-���`��B(���M豒�ܟ�"�Œ/r��/��i�䛓�*��U(�B @~k�@7�y	JZ�����h�',�����|��Ͽ}�6f�\��+�'��J� "�e����Y�T��Q�;�Fַ�%�7Шc�ϝ.l.�tZp�[������Om~q;q'ڟ�� ��v].����[>�/���1��J���O�qȌL��&3��J�vN��M �zBu��ח߶�C���7�ڵd؂����f�8�l]ƽ��Q�gPp)��Y������?ۀ�C<~>̿2/u�^��T����:`�o�)���'ΰW���UU;���<��f>nz|�u�]n�yHgIF��>,}k3cz�{M
�(et�c.iB�sx�d *���1�0�Ҟ±]�̊�U���(y����ǆ1憟��1;k��������� ����\���}���]��.�4�h�}?��C�3�09����L-�D�x��6��c��C̪[>�W:��� ��Tn�X�U��mI̮��ep�p���K��
������;��B�@6���)���$i}��jb�8U��݇�.3e��:]�z��4SH��$����F��X�9��33x8?w<�h��%��8��;%1��>{Ӆ������_��%�1�P����VW����iN0��Zϭ��9)�����\�Ga`�E�P:���.��ʲ؁�5��٢�r����o��Wmە������ﭦ��1ax��ꩉn�����!V����"�m����gC6�	�%~�/���,�X`��߱9����0�=��a�=3�pT��������YϞn��:W�dKep�.����Ը��#��7���jrG)PNL�j�X���?�u$((ޙ�͊s;��$�{�M�_b%lC�Z�*\����%�j%?�3��;�G�?&:�;�W���=[��Ϛ���q0a�ǲj�"{0��U���1O�I�9|q۰_���T��F��[��f�j6��~q�D,�_ތb�#fӍ	a�	��3���yq��[|�����C��y���i�1;�'�T�1y���<����%�~&s5���ټ�mgq�����Z�{_V3������R���Ir���P��d��%'t!b4RI��*jaE���U�PmO:�o�mb($��f�铍2�O���'O���?��r�E�u�DwYn�oY5�,lz�����T���W
����+Y���g��G�[.���9B��~jK�w����r���`���X�ץFw����j@�m�ďk*�`"ӈ�1�(n.3!��p�K��5y�Pa�Hq:�t��lߕa�*�����q�Z3�u=72	�Ε��(L>V��XЋ3�Z������HV����䅑��2��"Q�
O�������O�X*�2��Z�]��\�����` ��Iߌ3N��t�FCr��X(�UR���� "@�t0�G<��!(��=d���#1du�n]��԰�ޫ��6��r��[�a}0���9$yv�L����'x1
�]��ϊ�g�@��]� ?v:�Z���d���㚭~�i�+{"t�	�����(u��f�B_a�s9.�v˙�9�(ǖ����4�	G�q��,5��w+g��i��-��Lp�%&6H88� u�{��?��`����r���\���Ć<v>SM`��Q�d�"L�G�^N}��p��9��ȵs�/���`�UT��t~r~脨�,�׾Qz�7E��Ç�q�)t%��@l��3١�Xd9٦�ÈN��*�t6C�i���5[��l����<W	́\�Zk�1�r��H�`݂��@o�2�%-��'V�}"�;���!#�w�:1�B�椡vQLt�9��5��#����OG�5r�(��}��S�M�M��Q��y�wNr�w~]0ڼW4��M��O�6������5��L���@����#�hy�9��{���N%���Y9���Զ�?|.��+y�|�<�P~���5����;LD�V�p�<�T6��6��4��f��[u�Y�"�
�tB��3s�j�!<K�*�T��9�\�U��@������Q� z���Q.a