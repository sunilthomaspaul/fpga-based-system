XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��YB�NM�I��E8`vg��SH��
��_��q�T�9#d?޶tHmݡ�2t5���� �fb*`� ����t�QoL��=t��[W_�����a�N��┯�0/�wZJ����3�N1�����{U4Ss��I��Bc��n��K\��b! �%�Uq�4A�nMw���o�E��q���]��Dj��]��N��*zZ#&���D��Kt�S�>(!SNF��U|H�8]��Ss@�vH��^����Q����?��zk�V�g���[E�nՈ�Fg�/�k��*�Ŭ�� ��W�����6qPC��B~��?WE,bz�g`�5��밾�<����������O{��({]֝9N�|�F�BH�ʹ�۰�w�0�8��0"�� 򸻀d�&���i�Q�L{�9�X[�ס��qP5�yy�7�SO9�%����F��T1��|���h60]\�ש
�(]���B�mؘ���`B�
.��r�b!BV��.��t1��ˮ��Ͼjj�H$��,;���2�(nˊ^�XzF\��$&�tm�c}��,�� �?���i��F�5�Q�m֛������� �0�l�KY�ǡ��@_���F9׹�}7�]츲���,x���.����p�O�h��c�d�$��<�	�~���Ze�Zڙ2��6�/�9��JX�L�����E���t_����n�-\
fҬ�w�̙�X�\F�}�e��<yYR��1�O�!
��̻S&"R�����a�iX�İ��I/lXlxVHYEB    4c95    1190E�w�E�N��].��F^�R:{*4�R�^���"Y5�]� f�~DL�_��:!�xQ��gi���m`��}��9���_M\:ͷǱS*cFq`�;9�Svf�5�3���{�Vm����A�r =IH A��8]���>G�se�K(�{�'8����*���Q죉��-�鑫`���~r;�-�0���=8}oZMT�X{�����'��M �7R���_�E��~iP@��H:o�ƻ���k+1��іB}O�>�jo�l���Y:�F��4�6�ٵv��Q�� ��!{ʺQ0���`��j$34�(�@A�tތ<!�*��>�Ȟ��&�!e�u�J�QRq�V+��ik�UҔl�������D�CH��<.�+4�Վ��iV�B��m҉Al[e����V'�H������'	7���`��{&���U�a:&�=��_����1���7���`��%�����6���Я"@yfq�%����h����vƘ�) �ZpY-ʳC_;X�Z)Z�������0	.ܑ�.��*=�C�"�&�b�Ҁ�����P�q/����X���X����dZ�.����Z�'p�I,��� @����;��`�%���R�ֿ��'M�p�ӑ/���h/.H ƄG˘�V"MY��*.���a� Rg��ċ��-V�=�З��UV���CA�8��nX��6�ܖ�'gx ��X��@��n�·RBb�k�wwŝ�v�c�b�1�����	^����t]��W� ��΃��Y��6 �
���&c����^z��=�k�l;e���9�-MHơ>X�����C�&�����حS4�Rf���<�>v̖}�����t�5?.����$v�[��1Q`�n˳���í��@%���ͼ�x월�-���K�/��U�n[a��zp {Iž�RPi��8E�Q�o.e��a����Ca]@��|4�Dy�,l��f	Xǲd��]���
���Jr�:A���� ���2��k*oNN�Pj��u-���'�1.�kajB:qw���a(���@[;s�F�v��z*Hq�6�,}59�1,J��c8z�S�V��t��GXE*7���L�oуr;a�^��L�C�du^�vG��e,mp0k%�rr2\8Z��
��Y�൭-�k׹�f#�q�%$����CO�3B�*Q(*7�,��&q$�^r��*�Z���c|���Vw*�{�)7k)$�Ĝs��3x���ĳ��ɮ����a�f乿�M�?yX�eO_~L�!m���p B��#�%���uZ,�����g�g,1��f�Q���_,��j�Ð:�"W�SYl�C}���A�����y
��ԯ�R��w�qd5��¼��ޥ�'%����$72��\n�^��خ�[*�7�ม<#?j�=brw+N�����~"O=J[�s ,����f��������3�`���-t�9P!H�������Rf���X�B+��/���m�1��K��{b���T�.g��
�:M��5#7��ɠ~R#�'�J�.�#͹�ϔp�
d}]	��b�ߎ�-��KRM�Yj3 =(8��B��hU�����{�d;�^ K���T�~�)��/[�bX㦿�8�� ��*7��l=�@6�^���8��˸�P�<rzQo�艺lF9�qf�0��ADK���*B޲����*QbԈ�,��´Ȕe��=b��=����(�w�<��o�ǍK0w@W�e�o�>(��F$�T0�����ʺ��`��N�0N�giZLd�9�=�Td�Z�&	����B�F"!ϛ+lPa�|�D�����tռ]��"�~��ݙ���@3�e%�mx3
���&˿��r� -N�f���_*mQiq�M�pc�(�?�=�D]D�Q���Ծ��8v_�վ�ҔnO�U��e@�<���Z�q@*K�U��Ű��&)��ZÞ�kK���GAA�ov�c\D�"tf��Վ�7	@nZ�'�ϤJѪ� ����+͕�-�'�d2s{�ó���eXg0A8�@^6M�F�Jjg�U�2��ȯ���������D+�`������Z��=�� �UO���1��i/�})N�G����ݭ���\͓�3ڶ_�����_T	��`�mX�xZq����߆7?�&��0�nY��戌\���L�;F?�=��|*����8��m8�')���WvP�0N��)o�t����ܹ$:��N��A��νgwjo��9B8���1���}y�eg�����|�ĂK_�ڿ�t`-d��G��U�"nS�s}ѹ�����B��Sg^,�5�@�/��>��a���I^�0�Da�v{�'�z
�����8>&�u�������#����A�z�H��kz�y�
sH"*�ժ��}4�0��K9.ڰ����m0�Ɉ�B FW��ѳ`�CӜ��71Ae��0��c߳��=��<�3�´�T���ަ���%�ed��9D�s��v|�}&����q�_�8�s%R?yW���Ǿ��H�!X��6�/Q�8 �!����2���L��tX���]l��0����ՙ*��P���c�T��L[.��m@0!x�O%�t���� |c�cWp� ��N`�T��7V�Ґ.�vM5Ӏ�Ȥ1�
]>�� Ҷ�ڡ���=��+ p�4�ҏ&��Ǻvt��@ꯀ�|9/"�5��.����Ӕ�N��H.]eS=:/�Ky,#"����=�n�~:HI!��5s�Q��L�@��(�eN��� �F0�s�|v����7�׌�����	�������ĩt�T0R��h�J�I�W�Xc��k3Q|�1d�N�7����cۀƥ�CC����ՖX�4�r�-�ި��N_��6�WDH��X�����1�y�1�=����$�@��S�K�Hs�]�&+�����x��G�W�IX<�b�ΣY�R}2ڑ,����o!���\z�S?](��	IQUg���,,�Ni�s�$���%��_�g!�J�E��c��*�;͖ԕ�IPt��s�b
Pkp�z'O,X�~|{�;';ϊߜ/��~���m�������k�D��o��54F�3Ĭ��Z��}8�@=���!8q���'d�Sa��P���8��'��E�=��ra�N����C���[|P�u�?f�����F~ws`�� S\Zp>��@��v��A;iC;X���K.k簅��R�jO�?tk"�����36�<����h�2ד)iYEX(h�����%�"\l�ޤ���91N�6-�P~�66	hN�'��e8w���}Uj��Fc�&��5R�Aqx���j!�E�'��a��J>ϴUH| �&��h&�kZ�g�c�O~���qȓ9�8KӔ���!v�u�χ�MQ]Q�u�����\�	�+�3�����l&���3��yI�n1�>p�6��&ԑ&s�Or�8DeN!�� ���?�
��������J�K�\����3o�$�n�ل,?q�V��d�Tnw�>>���:�:6a��?��R���a��n�b7��ۻ<.Ѥ���R���U5}0�^F��F�|f�|��=�e��8��׽^�;�	%Ct �ܴ蕀Xׇr4P��V߱鑀na�7��s0��G� E!��w�T�,%��s�ѿ�ӛ�'@��]�0�0�����&�����ح��`h()�y܃uP�w�'4�=�Vx,n'1��K��UG� ��gun�*J�<)!�7PyoC~$h�3���0�4(}s�LX��A���3ڊ��q\Z�f_E �D���Ń>�̱����yp��7�L
�����&��c2#�Y_��F�t]�9��[6(���w��>�Û�'aO�̭����W�3	'����`K��{��磾��_E�s��?�(����d=j��g�Hv ��VF6���#�ԱG<��27k�g�2���D.��ܜtm�@��������j%�f��9�
oY�,��J�[�4K�\W�:-��k�+���Ll>�ui7COc3�M�L-�U���<�OI	v�a
�*�v!�2m��P�0҂0F��87� -̵FU��0U�'��[G�xA��ɺ��t$F���q5� �y_�@6�=e	�\��{*�:�}"O�����q��W��Q�Qw�����?�˃L�\F��V�!���'Y>AH�� q T��(�E ��c9�2f��!� qR���Y<m�ZjdG������j�ǘ'c�I735�6��Dz�T'�K!U
�g�q%��F3�5�|ɐ�R����-ةP8��vm������˴����*��k��t �/���K��A��x�f�u��s�4���"�X�)h	[�7[���
�4���D$�hW���%������]$�7o:\��/�AA5���p0\������2ʞ�
Ep���v����r�4�����7b��h���0̫-/���k�IT�