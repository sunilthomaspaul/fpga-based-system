XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��}3�M��bcȴ�ɧy����ʍ����{�jḺ��}�'�<����G��������ʽ���M��y$�'N5���<-(���L����ߗ,+�/�`1���.�u^u4t���B��m�U@JQ��ꞚԫT��4	E��ʽ�T�G}$��:����ZQ���;B�ﱕ�����mEp���Af[��'T��73��>�~>k����J�� �e���� �Vdr���*���,�ū������^��\<T��}o��nO̳#�R_�u�zW�{����-HD����j窀���aԺ�������3c<��ަm����:*2�
G	���d�����l#�!�G��ޮe����|
�N#�q9 a$'�/+P6��� X3��E�����S�ͫK�k��ǜB%�������{g���^��$�q���$�m�΢�7@�n̝���|�-�E?��:�r�]D�r�aa.�2��7�v�f�*ؑ_�^�������i���;�Q�p����d�Bc��U��9�.��6yc�7�y�[�?,O1@70�tfP�|�Z�/n�jL�Ct��W��ZT��Z���3�q�W�<o"�Bo�@�ݐ��3�&~�k/�[����$s�I[���ܕ�r�2x�����΄7-���)��3�T2���]�rZ��ڌ���܂����5Ζ�0�-Vz��cD1�ܘ������1�,�Q����x�T��i\v����3����P+-t�4�+XlxVHYEB    a19b    1f80������W�衵�4�,"T��Q�eyxuO��G��R����%���ۉ������OĬ�โ�A�,�bTL���j�͔*%���J�w�}ꖼ��o�V{1E���- PϷc`�&���s������z;o7RN��OIf��h�,��RG����H�����`�*tZ$�%��z���'$�Ȍ�����<d۠��7�^���!ۗoJ��$@(��5�v���u�x�#�,sx�SUk6q�-ǘ.���H�;�J�-fRJ K׿�QBh�U�V1�h��عۻ��x^P��,��:�>�$�dbI�������fp�
��k�z ������53+�7�P�0��8���A3�F���<�&�A�6e ���J:w,i�^6������e#T!�ao3���Le�E����TU���ع$v�xg�M�'ID�:gX#H�����	�z�y:�t�d��A��g����:�S�QGG�]�j�?Nqg���G.l(:���ZUK/��+�Q�r�}/�	��� ���.�P�}e͔�
I;-7�[|�����eO���~}M�u�I]E��u��`b�	�A�ז�0�(��V1��K#���f�ѧ*�"�T�����S�`AWJ��H��ğ7V���aiwh�ϢI�Nf��G�� �²h�v�O�Ƴ�x�!���_��+��ݴ��FF�f�i�����"��l*��n�5���/��L��?q��{�R1��\M%�!:Fq�;�48񫱬�c͊�Vs)rev��r��_��i6ܼQ6j��!������OϷ��8D��)0�����	�;?\@H���M�Y42�Z���y?\ D������I�u�G)y�ɞ	3�n1�Q�^Q�Y`O��PA�$&��u�o��g�й��Z2����Ί���t$�Z ښ!�_��)�ͧ�Ĉ�e*;|�B�e��*S�� �E����Wp�� � c�� N���/5�EB��U��SXY������0���G��&2�k��Sx<bIf�z��]�u
�8����P�+�^�pQ���l3sy�V�҉hK��?j>� ߇{�7E�r��'�y�Vd��P�+�/c�Wu+7��T���I���`ާ=�����z'&�<w/Ⅴ��!��k�)UD��z	E\��D�늜h0��.�혳"Y��g����d�l~���@��1�i�7�5��� �&�����4?��L���HN8����E)�2u�L6:P�gp�C(F�	e��28��5Ů�xΆ����cq��dѹ_j�{;�������'� �m�*
	�xLBNm�����t�a@#��<� ����
z2��
�-��\�a�O�J�gv��KR��@�h�X2�(��@�Q��Y8q�ҢYP�)���]�<����O	Ď�3f�d����̼7��~���E�'˛ۦ�!��Qp�)*���.ڤv#�H���HZX����l=$.�g/��e�ݻ(p_�ڇ���7�)oI٠���ߊ�^r/�/ϊ��2X�k��O[����o8ϳ�1�dIr9����Z�G��P^f��8X�U��Ի�$JEɣ�
�[�~�O��_���}Z�&�	 �a�XQ2L,�m.Y��#�"%����J��gA5	�z�|B��RU�/"H�u5�E!4���$'.�H3y�E��\J"��#�l�� nv��xfUO����t�t��PF~���p�p��ܟU\����>��O��i��BCSns�.���9�Jh3:�+�����6���h���>�A�fHR�� @�c�hp�8M �*V?�,�V���]<����$? >U���bn�`)+i���ˢ�Y>�7�YJ.��-��F���[���+���*dz(nM�WC5�Q��J�2�m���(io~�v�9
58���m¯_`G�%�Ʀz%_%d��#���P<��䃳KQ�`��I�DH������e`�у9C����
Ք�h,�#-�_@��V�+wɟ��p<��.��7�r��.�t�:IgI���J������4�p������v��՝)B�`H���U�1h�r��1�%`����W��y�l�ֈ��� �J��F,|�_����4Ԯ��V��kΡ	'��k�;3O�2a�Y�s �[}�A�[y>	������PR��$�IՍ-��A;���K�r����{m2�?�:i�h�w��[�˸/Aד��x0���.�����ْ��ͽu��@��|2�/�;��m��B�D�ȗ�D=<2������#Y��BoF�'M�@�zcQ�\'i�?��ENx�"��K@}6�L�'�l\b�3X��FO��c[��DU������Ux��Ņ��&����=����Q��78�0%������;�ZC5c�F��b�S1�z�#'sK��;���7ũ�\���@�6�Q����D'K�Y1����#,�o��{$�z{��7�fM�r�앦�g⨆m�b��J�i�P��8	p?"X��v���NC���iҺoׂz5��:������k3�}h�<w|�]�6d�%���I��դ��g-�d>�&���a���x�R�I�*�|휦F��d�%0�xw�7�:��8�^�M�2�������ףoX��/7$r���E�����&��$�<��l�{��
�jE0��䂛�%x�{�M{�g�-����ރ�,t�b�s)ON_�Fq��m�|w�"�.P����
�y��ɴ0��$����nޖ�/��`H{C	���V�d��Vp�尐�7"F�B��#m�m͚�6����|�"� � ���ZM�@T����Sp��$�j1�=Z�$N7��.�.5b�A�7  I�$�֖سy��+���G��D>�����P#Q���C�}�4.U�N��W1��<N�*-�4qlD?&��t��E�G�����"_�H��u$��6�q�n�I<+�y<����/�%����}A@���������볚�o�2in/���k�f�oQrӇ���/,+�Ê��m��ےd��o�)a��nνb$�d�Y�cO]6=�H�*б�E�r�	�ƾZ4�N�fy�Yb�5�٢R�y}��HlD	rѿ�oV���Z[N� uT� i��(���_�FA�b�*A06�)����%����?o%^���"�e���+�+dE>AB] \���,��}T���I�$aI�hg�Ix���]L�����
����Z�O�,9�7⢟PT�������c�9hq���<��4����<;7����Rv���,6����XW�i)V��>���q�����c:��S�������c�(���	�j��l3�>u(YTy�ݑ�m�] ��=KU��>���[�uR��@�Ӑ���0ت9o�������[@��!�<Kt��G|	���G��Q���=�[��>c �]N�Oq9^�n_���1;Kb�wS�0��p`���==��NjSi,�� � �:���`el!��>9˱U�G��F��ѽ�:������2[	$,��2F��(��$�"����+l��3t�5�!�b^P+xDvB�8��'���Q����dQ�L��Ve���W���ӳ7�c�VBhq����%����C�`X	?)���d5-�tT�_��r��,�S�`���/�M_	�,�ϯ�����o����N���u�7�$x��y,K��]Q������	Jq�E5��"����_���Q���=���T"fVr{Ą۫4q���`II��	�|$y[[æg[Ԣ�6Ҕ�F�2�p;TL��d�VS�}�+0TT�3_[���"`%��Hh�h�����l����ی�PT�g�Ѡ'���:*��Ȇ��h^��	}u�֞!8+�gD��Qoq��Bd�RM�ѕ����ؾUz��ʋ��È˪H�Q�"�Us�gψ�!�OkH��U7V���Ւ�≋��}��5W���{A�#ۦ֗p��@fR�)Mׄ�%�l�-:��ʘy�I�.="IA�y�l��n�$��,���9���-+L{��(�G���u�v,��9[BH�y�����Zd6�?�!�8��������_��ئ�%M:�cz�BI쬵6�;XF�.I�V ���g,�e�
�e���>R�G4v�Ϻ@$��5�8�%�a�d6���n,1C�����ԭ��&E�xQ|��Ӹ�kM|P��8������#���p��)���������9��A���ՈߛT����Ji&��7��@�z�� f(`]?���^5L/Zt�&x�)�i�S���]�2�7��b��{mt#�;��}��w��U����SA
^������|3�#����g\�FPbi:uK!�Rw�m;� k*�®�u=�ʩ��*0��r�  ��@�*�4uOC���b	9P���k��:Z�{��2݁�� '��i������1h��|^'�m�[V=,�_^6F����pT{����w�ڜ��!��kPa� �p@��ρ�Z�J c8*�.�|n�AU�^ƙ��,�'#������9���v7�2���E�@�~�47l���񒖯�ݎ�L�2LJ��枒4\����U��j�'I�l��*���落��ɆAL��-�W�|dn�"b	5q���Jr���!���ϖYyp�v��S�l�	ƞ7atMG�����w��YT�^�^��!;�C��ʩ8�|� �vR:��%�xf8��C�_��C3�7��/�_sD�fߴ�j!�.P,"�=t�%�Vi��N��C��ʦ�)s���d"��H�/ƀ&n}���Ub�X-!��� ��I�ӎBP���G��1x>�8��L�%o��|<HV<���
#�ˆ�Qǧ���\
<�Մ���K��cZ�wA���V����W��f)�q�%��8��r$ۗ�䗧��9*DU����2����T���7��0h��9=Uя��ϊ�{Q�=j��<�i���R<ި��_��{
z{+�
�x�4��֛�@i`6� �(��Y�d?�;�c�o-�
z�;�X��"��dS �O��Y���մ�?�Y7�jd�Ţ�*���J���ޙzЦɤ��R�,�10h�`��bX�YC
1�JR(�a����b�o�i�Rsfˉ9��Ǯ"���tH8 XF�.д-��\�;$�Q�iJ7�(�(�!�lv�ܵhk��y �͇)�Nt�� ISZ����T�{�:$��
*R��kTU�����D/�j�L�@r�I�h��f�]%��:??�	��>�g�����P���xE��QY�F҃W�)�U|�<�fK�5��t4տm4� D��3=L����޾��&W_��2��4��]��t�J��	p�Po
[��O��m��nJ�Xe�W�'d�_���]��Xes߸���og���$���)e֝y��A�OFd�E\L^D(�p��NiYjn�7��@�J�]�����2=m}���8��������-���|��ڢ�P��)f��v(.�%^���5�;�Nt��)���q�w*����j��R�Y��w���KF_�hX�{�$8k�j�.��Cd�/<���e�	�>Wl�ޓ�߹��4m�?T�$����S6�W�$�=���F���cM	Ӂ�dM���؆ڀ�D����v��WU�o�"��n-Y;jY|c�tf�%��0��1�̿�ȥ6��L�ө�c����0J����~+Fu-�p�h2�8E\���_��ړ�4jﵻ�[T%�� ���.���^x!3Ai�f���.hoD�@��84�0�Rh�R�B�i��´V��]`8�S�	n- ��3*��zگ��pk�6��s%myQ�SWu�@�ڮ�nqgꎠz38�S��'�b��n�~+��F2�t�U��i��\_�B`J�%�j��1�"�:t���q�M0~�ӹ�9B��$�g�S�4x��w�l�ȕ�������x��r�6O�˩������?}�Àȹ�M�	���i�$�Ԁ�6��0�D>k���:����u�qecʐ��\d�x9E�[�+��}�c�_�(/�����sNw�un�0��:,`�y(���Z���C!�Pk;N_�[GIB�Pa��EY�J-�?\<X��t-��v��-���ʾ��&%u���:�"��x������%pk�������A�C�+u٫V�E���o$�Ae����Q�3���`�.�]���$�ҶՔh^�|�yv6rh��q�Q�Zdk[s�<��<6=����~���^��T|
A^E�b��]x[@�5����.�W��^��uU�"r���0�'�������p,�K��x�Z���4�5��T��ݜ[ς�v���r�:}w�UT##�V,7��q�%	��~y&�o��c�����y��v�����R}���W��Cf��������M>7�_ ���|���t]������2'�O���B@�g�阔a#f�f8�笪��F�N,VA>2	 .�g�[��h��%������0u\Ű���ue
�-Ąj�kɌ7�5��Gsz���[,��#�?�_q�l"�jV��L?���d��V�O@N��Z��0t�s��޴��4&8���^&�k;��%�V���W����I{W�R�����&ԭTQ ����<�#gw�f3�t},���/�TU���Ď@
�(���d	�+��h�j��]5!za.z?8��\s<�Rb�SY�U�G_�/�4�#x�b+v���|N��]<״Sl�m����`d�h��P�{�Xg�u)��6+K+�����D��Ⱦf�Ҧ�Xi�������%˵�r  0ůi�Ko�L���C���ؓJ�N�MŻ��a�D 
\�?�Xu_L�ժ���m�1�K�O'B�zo�9�s�w���RJaW�Flp$�ҩ������vѱ:Z..}7T��Ѩ+X%�I��W��r̅����\����&�.�P�89E)��~!g�TFs+W�+�&����8v ͬ�"��Z�CZ��ؼA������KV6}����8���9��G$DҊ��pS�Ai�<ѩ�C����:#���""Ki���u��֟6o9~N���%�x�B��eZi�1�0	Q�lq��o�nv�cG)�T���x2,��%��t/7�؝�2��0J���I_�53����})\A�]�-�^���+Zp>E�D���"�T���!E�G��R���=�z��8R���d�92{�0%�ܽ��@,$�\��c�驭t�N�]�G�"E�|�B�C�e� 4OGP����I6�5K�U��+�?�����B�Q5�uOS���`g,���7@A�(V��ca�0���S��D-�;�߫�g�-v+�J1�ϯ���t�y�Z������9����3�����<e�O L�� @#��?Ϳx�0rS~Waʩ��lQ҈ M����I�q'�J��ȯ�r��5k2^��lH,���jP>8�zky���%N��.��#�N�a[_����>q�^��*���_�.�0R�`�^b"M��#��� �؋	����K��L�䨋�,����!�6�:�Z� m���=�2�f��al��R��u�Е�>?���0�g2����m߄���1�=� x~oz�H�=����6�4��Xo��v��A��~���{���N��q~Ug���Θ��-��M��i.I��
��-��M6N�rIL��Ħ[7�{u>���A�iS��K�<^<����������u���$V��Q�F���jg�~a� ��Z*W�my��[�z����&����f,�u����UA6%�U�s#�`r��:t���]���ˡeȮ?�Ѓ�__��L�8 ����a�v�f΁� ����=���K����9�_��N���)�iLc�/�-�x�0��"���ǶVl��8�%�l/�fG�9*�:H��J�H