XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��U�/����h~x�]n�݆��2U��^ɵQ�y�|�ڍÇS��@�x(<���ss! ΰ�«r��+={TS�u��,G�Q�t�3�FΊs����2^�в�<)������@�!��14��aA"�c�z̆#���9t�F���|5�/\8�0����W���d�����Y~x翎���EY���`\��ܲe��1���?�m�U]���jc�f�IM���1�YcK��XGH�<GO���%s*X���S���'�X�J3/q�{t>]���Y��͔x�pm�U�߂�.+����v�ۅ٘� pBZ��
��P��g�	�A9�Tr9�z"O�����w��"��΍5}�)u�M����U����ep�ી�M��fk
%�7a�}q�0��#�KR��y�1�H7���]*kr�И�"����)�ȶ��ĺ���bu�,W��Wl��`?@�-�8�ш�3�{Dw�+?EuY  s�QT�I��]��r�c)�	jC���ȷ��N2]�偵�ʸǆ�7!R
�+�  ��>����x#R�5��Cn���q� �z�7�?�&!.�!9�Zܱ/U�V�`�X�W���"���T�;�{��b�}c�)��<���/�>� �� �ތ'4_j�U�+�݂��Q2fљ_��-j����/Qo;	��F֕^s�օޚdrQ�&������t�r�[K<�i�>4��n��/��0�	V\&�q��;H&k¹N����-�XlxVHYEB    a19b    1f80U�ZU9� 8*�R�ڇ��i���gz\�D��2�]��4��bY"�^�Z��ޝ]�z>��o�d��߅m��OZ�'���hT���NC��pCV�_�m�ֈI�����U7ؕ4�y��a�9	�A�������%(uf��"�y,��^A� q�եY7Է�0�.6E
���U�� �����  &3�ȥ\܊�׼��1��b������'O67~(��Զ�Bƫ81m�izK�5{O�t�n�O�
*aY�]/i��'�������I3W\[f'0>NWDDu��n"�ƴ��cƢ9;N&"�טӮ��v����*�w��Q6{
U��Y�0N���3�iz88lN\����U.Π��N�8�knU����Qҹ�9�ω���w7Pa|�-�'��m�C��ٌ�r�?�Ь4����TlB������S4F����N�y�Z�|5`iD�JS�
]%�J�`v�.8�T�AT>�������f��|ŷ«���Js�F�;U�A����E��?ّ�ɾ�B�1i�ul���ai�"���p_���:/F�h�uW�}r�h���ڐs[��E$�ԛPW3�~��_t��GHjp��<C����c���Ȭ�K���)d��DE9Z�+��%0����=����U�\y�����Z,O�=��c	�s�V���֫.Q>�'�lR�ĄƖv�%K����F�ǅt�Utu��q���Ⱥ��o{,����ڿ���N�U��y���XȡI����� ���LP�	pO۷;�S�/�@���#���o�j�?��n���a�����sL�ËH�t���th��{�c�9RU�f��U,$��y��a�����Ý�a�aq�.s�ө�װ��#Z�������\%!I�ED����G�*�?ن
rz�/G��cq'k��|����F�H�6�Uks���εg2�Y�=d�75�M���3H�������nW���{��j�vǑUA�.,����=��E.e�fJ����f��ݾ�Am��8����)�qb���3,�q�{/����+��ǉ~�bբ9�W���Oitj���sʏ�9����_��
#�O���JQ'F���J&�� Eʸ|��36��U���g����{{��C7_��E4�R�lx�)b��Ũ	O"����ݑU��G<I�:�f3��u6���ܒ^k#:B���2Rxk�Ct���Y��˔�yD�����H�m9����L�>�e2���v^˔37��i��@�0M[��}��MT�T��c��Q�X�]y��d ���R%�1��K�aj!�f��4���:�̤N-�5vg��C\���g:F���#G�V$7���[b�9iR{{�Ǝ��Nn��Ñ<��T���¦���m��R)��e��Щ�+�ľ�86�Z-kB"��W$���L��ӥ�bu���T�)�3�K���<�4�>]w�^ܛK'���[�Cƈ	�	0�(���\z����z.�?�kKlAk`\�^��َKD �Bg�/���'J(B�Q�/��B�OBdҘ��5s+�4�<�>�<��0O�@�.PŜK��#�F_&o��8��s]�Y�C�86}Ǫ�e��]}KD*����4w�_�vAF[t�=�(H��g��2t�z8N��_��x>���֘�jE ]�J4J�&��ÖИ��I�����f�N�P��my��_��^~�T�C,�A�T���;?�غS�)u9�x7���R��=���_�u��f�� �;49��GhhG�_����l���|p��A�T|�,�)Ca�	0a#��x�<`5�>?�e�F���i�����Z]a��H���Ԛ��p�t_� �zn{KD��r�o'�ml�uEw�ɇl�x�:�	60�����C���Uz��M�X��!����]�c�4cq7;����y���*��i�θ<
Q����rG���ң�[B`J�D%�7��+���[P:�a��iZ�zgC����"�
2M��e�(;�7o���$-���<j#�q��&r�����V��i�.�Q[�M��x���33���/���s?�m����m�̪�[@I��j��.k�U�$��0�{�:L|�A��H��'!�ǰ$E�KN	��(��z��^T����o��+ɇ�(�BEs�+�ކ�hy�>���6 W�����K�v�.*�JfN�����/˥J]r���I�H�UȐl�wX:��#��X;���ӆ��r7����6��(m3T���7���V�-��t�7ؑ�?��#�5^:Uz�.=���f���ga�w5��w"\l0���hVެ@��*ϫ��G2Iab!/o�Q!n�(؛ݶ������a���2�+7����!�?�ʇl�HWυ��*�'	�%�v�C_��;��(��#��ԛ_��T�%tVM���4҇��@W����nh��~�$���q��FI�#�[*���t�����v��-Bh0����й��O�bTb;_��k����j±����G1�I  ����[��*>��xH�r�:6�J�A�wF������+�u�����8M�r%=}/�Z�7Q��� Kd$#����,��� ���fĂ�����v7|���UjgV��>�P��������	5�$a�Ő����ґ�u!7�����Z&�~C�L�K�O�k>�����n���B�Y��׹��̈́���m���t��y�}���VV���HK�?�[3�_j�	镱,};�BY�`�K��V�mD`]RnX�5�*�.3�5<�>�J$�V��>�buw�X�At�b.��ؼ1�\��&�\��#Ї�"���7��;�\�ݓ�{�N�F@$���DYg�	 K�)�7-��� ����Β��pw�S稆焭ǂN5�Q���f��;)�{p{����/��H�êԅ�v�=o[膲�J��F�+n`7r#bu~�8�_(X��QE{:�r�ۄ[���M:t&���p���Ĺ���x���s��2���_I��]h�;�0$��"��\��<�⸿�IX�V��/%8y})dA��g���=���K|1�� �B�o0G0�qS##�?j� �bkpC���xj�@�I/ʜ����q�����y!�������um-�����.4EH����~I
tUB:V��t��,���!��7�m#�	� #��$j��t�a��H؍��ݑU�����9�K{��ٱp�-��Mn�]��*���� �9��Yh��<����oVA�CK�鷗�4vUL��'�~��`J�V�4 ����+���z�?�Β�[y�~>w�M<Δ�n"M^�]Q�c�eb�_�Q����t[��%!�Q���JM�F��ƔH��%�&'}�����N˜�kJ��@0b~a08�e�ZG���	��8�KT�	��C�i� �$4y�U��*(qU��g������|}�`�R&>���q��9�>U��vzX:����3)Hl[_����֐A�z�a��>�9�A���#Od2�=9 |֒r�pS ��!�4l����m$��dJ�1��� 걃����c7K�'ήS
��� ܦ̻
�B)4����)�5�/o�1�i�4?�݋|Z�b�b�4�����FH�+b�a�!�V2
�9	c��_���A��7�a���|�>)�;[��F�ou���w���1i̜�6WU��H��dƨ0N.��(���n�ꠔ>l���P����A	k33�ׄ���$��-1
��IZ&���k��4eLƂ�����*��1��P�-��.�&*�k�4��<���p�B82ӥ�j]~!��8����^�Fgj�~�Z�a��SQ(��GB�HĔÄl؄���B��I�r�W�o��]��%��W�JEQ��CQ��H�zh��(*eZE��+rN ��aB�8'�w���y���m�}*^�T�~���45P&�F_ �i%��c�[Vb3�f�ˡ��H͐�R��u����Cz�X��%��驾���=3��5̻���(�B^�c-�$&Ѭ�p�S.#q�ѽ�	G���*�Ա1���N�Za�8���9o����Y$c6�ܝ�m�4��Ru0��ؽ�0�%��7�<
�(����2t���C��SL�r&!�3q�5sR��˯��8�Bk6������$�L�$�_�ч!-��ʫSR�|-Rm��{c�U6/_X���M�>���V����{��OB?4��O0(������)PD5��t���z�c骉�/"��U�z��eݵ ������bϘ7��,m�O�A".|^���ol�h�?,�p����i���t��9�"�N��V��z�4{��ʰg�ۇ��۸^�V��VB[;��L�}��Ks�ŉZdgƱ�o�+rAU��1)b<�c��N�0���Jl#�{�S8~/�t_V�z���@�6���) ��hM�l��}cY29/Ҭl>�}����<j�R§�L���E5mJ�(>"މHa�O~I"��sE"Lcw�:ȋ$_��r�c���x{F��dd�ʂ������ɁHmQ~�������خA��0�(#|��*c,v���x�qT��6(T~@Q�����e�H\��9X��5C�'�4����D�A�C��l���9̛%Br�B��kZ�$��P}����T�?���~=�a.7��	�,��	�j�9�[��`�� �x�&��wF�i���'[5jbq��r�M�W
3|��^˖���B������Y ��^�'p�I����0����c��$��x��d��_0|Tɼw2�rB�F��w�/?��,��%|$ �s���e�|�d
�y��J�Me6g
�W$G�C_}��>��� �{�����}�n��T ��0H���g�.F���3�!��Ɇo�(i�T�����k
���y�$s�r���v�|���~��><c9-�|����ڪ
:��������/��f�����U�c�к��w<�����:�
��ʯlB)��!Y�B�����W�a�����D��~���3��`�\(&��G������w�!j�f�ˌ5���ܱlo����)�t���yŚ$����=G{�)���p��$a�KZ��RF�}�)���M��_�����hh^�y�L�(��D,��HB*7C ����Ьfe��{�K�F�0��#��<�Q�S|J҆�'�%Ʊ�}�(D�܅8�ޥi&*��E��Yg���'c�:u���U�?�5i{W�-��	���F�t�<��\������+_�C���5k$	*>��˂G��-�H&|F�4���+�����㾥:�M�eٛ���s&�4Qa�@��,�i^ia2,b��ٺ'����
�����M�i�ÊB��3.�@�X��W�V��Q�d��$���o���=����2r"�����s1q�A|����Y	��i.kS*�&������S�J��IB}�,��O�L�����i mK�ȅB��S�x���&��©�1.[F� EW�+B���Y_����0�,e�n7ʷ��R+��G���/�Ћ��ϡO)?#�5�ҿ�� ���FE-��V���8�G��n�vƓp����I`��|f�W�s iw]m��S'H�a<Ѐ&�l+��I'������K�p����2ӕ�F-л@�-�D;JڮIos*�(�D��V
򎞡>��U�.�/���q+`��f������?��q�=s�ĺQ��h�|�N8(�Xզ��%����<����!l%�J��JM�ܦ
0��vc�.mZ�%bڭ�.�l�y+-v�c\�/��Bgn�˵�ѡ�$�n�2��޲G�y����)(#��gg�h����&��Z���ch��Q�v�P��'�ѲA����x��5����L{���%�\ܠy`�|�*�S�y��jRIG}�}�1���Nu�/��%bu�VZ ϯW�a_�Cy��?��0��r�Wu�n�s%=��+d����cH?`��̗�&|�1M(�)���#9�$1��X+A夠1��-�z$��ܭ�MaQƪZff�c�6zٵ�^j>3�w=˄P!��G�X�aNJZ/cu^�Ol5U�j����%��2"<�V��{��;N�Q*}��G�c�d_s�ͮI&	>
�v~�����ۀ8���W���n�!�vKP*��2Nν�T>(�LX֓���x`�� 7��N�m�� ^������.�5��G~!Ma�C�Li��V���� Q��I�9wﾞ�"Ϭ'��F� �� 9�CS�,�+�Ժj#���za�ŲsED�����{�p�r72�s.)��{:�md5�sHؕ9��&�����?�\�����r�s��c���x�lv(�&AK6:вz��3��r'��æf��g��8��8�<9��rP$w�a�p�ގ�����]2��bYkޓ�f�^pwH`��cIo��b~�:vX�]ܮ6�	��J���$}�ٰ�T8��h���Q�q� �A��?	0���
�t~���АW���,εH�lx�ޅ�'W'��45�|ڟ�9w����w��٩;Ky4�	d�P��x���n��N��C���������)iP,Ⲥr󏢑�e�@�U�u%�N�*݀:]^�&<s�Hu�4�YP�Z�kW���ߌ����=�S7ds�>iE�c��ǫ�h I:n^��%3�0J� c�=�O�-A�.Х@
nIE��-�L�2N���L�NR�n���� پ��g�؁�����P����D)g�o�S���X��e�<
����a/��p�kh�c(dl[ҶOt|��3.6!�6�e�	�W��F�t��^�·Y'j�6cU"�ά���F6����H��UW�3a�e=Q��ۭG�,�q'���H�����o0%��R�g���3�V�V���Aډ��Ǒ��Q��]d�N~�g��]��/BBx��Ť�,͌�~L�|��@��8��޷G��#�s����Q�+�vXG�,K
��9����X~/���f-�J�%����9�مX,d�7�I�_GNP��;<��!����G�q�ӟ���{�~�#��bW%��r<�<�����1�m�=X5nG�0�/3�=����#BL�*��g��D�S�KP��*C�喷��;F��q��@EZ��4֗Ek���]R��l*��D<�-Y�H1y�-����' �;~yfa=2�6�[t�N�=�2�L��'f�����/c�|���e�P�ϟG�n���C�rףR.cсZH%��&͊t�׵�J1�$N�ġ�00Au�Vm� ؐ-������-_5/�ӫ�A�a2'4�����($�~���2G�5�,=NG��H�@�SB"r0�o���S����g�&�©y��P��<ꢥt�̸%�+9�Ԥ
��v������/e!�ӿ�şE��!�Y�0�Ȩ*h��
��YTlx ?��.S�ڋ�Zy��Ǣ����;��}o;��V�<�Q�:%��������Ŕ���Τ�Zp�5�T������'����!:>�����`�Dqم����K��k�d[��Y�0)x���6H/#l���:>d�K��lSnJ�Rhu״|��7b���a#���7�$C)�Y��2�����d���s*�o{WE��8���ܽTF�uJ����Ҭ�9�����ef�6~�8������Qb9_aB�?R�}��}�ˬ���t�%/�M`pʈYҮ䡚����Z��V���sa��w*8M�Į�L ��x�MAD��O�d��m�}\��=��'<���%~����n��R�%!�.�#�UL���׍K���������ѱq���g�	z*1����+�b��y��v��y�J��p���KZ�Q�/R�Ϡ�6��sĴ���Я��Zk�l�yV4���E�D��E�xK��V���Pl��W �୙|S?'\���t��A���|��i8O