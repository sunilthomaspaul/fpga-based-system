XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����H�M��啉q����O��'P�� g�<ԉ������q�t�xm��S|vd����Su.-Tz��#�!(�_�̯���$}��:ɥ�K�P�>��ɠUJ�UW[��o%q��4��8�`P��q����qs��m��A�M���� (��e@V���t����B�+`қ�QȾ��pj��D2��D��ג'7.����K����+Cddt�!�O|�Я��5���l�u841�4�5�V�R&F����.=�>_�Uov�:�����$��]�a��M����(e��9��)&/.���(�XW�D�麫�?���D��0���nb΂��=�{�'�9�B��L�O�*�,���Qr�`�n�e��qN/y�y���1"w6���a�kSa�7eݻ켐B|��yu�E�t鷏�9B�o~��Rn�B�PT�tu{`�3d�Z���n9�����>�ET4=%��|z��I�w�1�MB�N7g������@�*��F���Z,���q��(�Y�-�e��/{K��hx=���%��)��3�Q���-=���e����_�KR7=_Z���&]��{7:��n݋f�%�}cLR*�����R���j�����D�#V���[�D�r��}����->�"�!
o�R�1-��߂�� �E=����s&$�J7Ք��I��1��g���r<�^�TW~Bܕ��C�a)Wj���1<��b"�ugU9���7���~��ͩ��ޭ1!T�GT(g���(&���u�>N"XlxVHYEB    3e0e    1150WX��5g����y,	Q�:����~^��4�!���Ǎ`�ւ�7Q@2ޖ��F�0BE���0������b%k�N����H��y�R�0t�0
�@�!XT���U���0K}ÉHCo����sK#�����V+U����ۂ�3��Hy�vn)Ce�F��n�!vԁ�CIf_WHՕ�s(�.�$��W�(��@(��̉y��1��-��DҊ����.�	����u�u�n�d
gR:�1��s��?�7��a<���Y�C�"�*lK쏳/���)�+LcC�8�g	o�C�~q��p���&���蘢Ru�>��^�c�0�C�ٔu`P�D#|YQ�@X����y�D�D2k�X�.޴OMVO�L�k��1󥰯L��ׇ�lC��A](
S�o���B�����%^�
�������������d>@��o��jX0�X���`��y�g���`nk:ߌvx���p�9d$��g�qe硞��8�OP.䵀�&{|�;��%�Uy��X�O�B��4��AF�z�ÜJv���������,:m7x5R*G�)3�y���K�u��2.�]x r����B�#jȍ� 5�\U�4؍����%V�ͥ�8{O���f��d�d2������Ǌc<Rs���� �?��ݺ�X�M��D5��D^��(}RߕG`���M��e�O��nZqB�ň��������-U����0�6��ClgyE�\+�4$ ���iF?X�U�E�W]������ 7����E([ۏy��.N�:�f�#Dh	��Ӄt�������B�/?}������|�R�'b�<h+U�9�����[��p����.)`��	��]Z:(8$
1o��2)A�=h/&h
��9|>o�>r�s��|� �l�q�F�U�6B�Q<ΥZ�&M׋~��IG�(�U���Q�B�\M��}}۱�d�Ә�%	:7�(4<�����o��]�����B�`�2����Ψ�Dd3�N�3�s��z[�F1̸X�ud=�>1:<Kx�b�%�*��pI�'"+XLҡ �U�_p�P�w�C�����G!�^D]W9ٞ���|�RS����#�F�D�[�k�8�|;=�μ$�r���z����x[|�����?���^/t�aKD��Pp�IԞ��5�dv�Q�:�Ļ����;�-׆�#V���g�<Lr�#9�Q��� 7���|����KҞ2�$�q�Hd��u�nC�@��ƞ�o,D*��b�ᢀ�����ش��RL13UL�/5�t�5Fs � _��$�o���s��T��"�q�j����^��}�j��"���w;ܙ�����#g�-�Q�3ns]P���&��V�l��������ӟWI4��,x�%�~ټL�+���[�����0q?�z:�bM�����Hx�����2��v�T���ɕ�n(��q���[*��ٛuDҊ�s�E4D
<hI�'�Uմ���ge�,�+e��E�&��m�i/`ո/
�5]=#b� ,3���o5x�2(�C��[�������_O�M��"*@K�������L��7I�V�']��'���v	�F�HH|G��gKr�%[�G�8e��	�IEoBejy^��YDdw�g��P��C�a)�C�K�J�{R"=���Z�f�P��m�J��qgƢ㣸���^��!X�؉؋gǊ�<��Iʊ�հ,J�B:L��	+��|�n ;�[#�C�|ɵ�+�U����Y��ƶ���_d2ڪ@cv����]�^��4l� �)5/C�P���?ok�M�Ǿ� =��U>hbi��t��n���u�B5�9a:q#��t��$M4mBz�B�Ԇ��6��1$�aNw�o�d�}�_o'Z�2�Y�0��m�������/�0wz|��h�uYs��FWM;�����w�6�r��jgDɌ�P#+�/���H��� %�5ڗ,��d��^��}�m��89�;����M��*���ZfC��b;�H!�s)`�?�E&��:�I$k[�ܝ���$7g7�����Uu����>���t�8�e	����F����t>2x5�i��ʤH��������f��sC�z%;����xrFh�V����(����ep�y���]�b&�4�1��[�7x��J +�M]����c��'~�ë�`��q��x��NH��srvSar �. %�Hx����s�$M,k��sr�-��-�3�bJߩ%��FY>�yFT��������~�7�s%�o.�m�D��}�x���[��F�t�V��iZ�:NSH6,x�P�E]*&A�Q�Z��.\]&���a��t��?��yʶ	�I5~�^���)!�������%�=�(y��)^�Xc���rȀ��`I�B��-��B�^�W�6��x�`�W�n�Nd�eL�I��
��X��<�Ԥ8� ,��y���܈jH�"CF���pkܪ�ě�k�y>���~�n�z�I�&�h�ěᲃx�\��O@fz�a�RE#'++��3|����a��{��|�7��m� =_�
,�Ի��=N��FX�j2�W�aQ.69�|�4ݼjF��*yl�m��8���7l���?Y����=�1�����Hƛ��D�ѻ���p�ۗ���
����;#g"l���Ʊ�׶���2:��e�N`�{�|@Pᒟ/8	pv�_#�(nҏ�^(���H �>��	j���R3�Ӽ��DRg�i�-�^̶�T��4�Ĝ�^���p�Ӡ1jCk<q�Ϋ
����u�RI����R-BSWB�f#kIi��)�ꏠ����޾��R�n��B;ŏ�����5�zGUQ����\gp�79�Q\
1J%
�$v;���>������3\N���09�%~��a�����5�m���x1����bݟ�m@Oq���� :J)���z1`R۰�ʋ����*]���������!� �.z���(�[d�q�n���b!:Ϭ*���f�7C y�!�Q��
�OHX2D�����'��?S��zNJK�|1OB�K;��=�uD(0�m��N�7U��T `"�պ�kWo7������:�`��k)�f�!��G��qX�6&�����-��*��^�(T3!ڌ^��Q%6�*�;���Zɑq������f�x�t��೭�w���|_��}PZ��'r6d�L�[Z�\,��E7����0"��I��j1�C�!�z��_+8�B��Q��b�f?Ϙ�4�� ������x��9�3m��s��kW�{��veRfl��g˕�退z`�JKnX��i@2��('^��=/��޷x��L	;��Ӑ��o��}��旟�����k��ޡ�}�]l�q�I����:D����f�����$�~�� E��<�,mV�Ԃ��J��Wќ
M>�Y=�b�/s��
K�=�����Z<�&_c��/ M 	$�)&B�<��e>^�d����
�	��dM�Z�J)F>�}�X��:$�#��H��Ⱦ�q1���Jo��G� |��$8�ɴ;"3���h����j�^�@��{-ѪrL^2�GG5@F�~�-�|�=�7�y�Kh�hﮒ��P���Bc <�n�v3[�OM�n�.p�m����Y;e�ȓ;;���no[.�H:J(�������^�7�p	��-`�ùe��]8XU�v;}W�F��-W��T�P/�z�������)5���ӱ������I���ys���Nӹs���� 'H�K�T�ƶ��zO@�uQ}�*����c�99z�&�h�foV�k??f! IWax���"�
����՘��_�}������Ң�[����������H/��k�j��u�z���1 �+���� ��%��l��J�6���>�{"2�TO.�V�h �~���<'3�	��J@6E�&�A��F�L:�B�|b�#�\_Z���k�VOA�~{
FfL�nE�L�t,��G�g�U���w��D�P�Իn�$�� k�*/��ޝ|,��\-U�'�����D�ԟj��{�q��3?���J^����30īO&0mw��[�S���s�DG�*�*�<�#��@���r�]@�e9pY�F*g]�͊3c䒶W����^�  \���׏��q��E�>Ko̿����9�v֔D�J4kwف��&����:u��>�˳z�i �e{2���WY	�Rgle�i'U���o)����v�'+B��J�@V|T�v�ށ�Tq�6Qm��?N'`������=��i.Y�.r&V%]�60�#�V1U�=z�YKGr���5�g��n4i)YAo��1B�P��W��0I��W6FC*�wd�p��Ű