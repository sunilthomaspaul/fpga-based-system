XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����w�@~��6;DElx�^�zO2}���`Ӱ93l�wum}i��\�Tɨ�>K�[�ֵac����:W��5��� ���!De��r�U����]h"/7��Miۚ�� ��|�P��l���f�t�W��z\���H���l��|������;�s>���ϰ	Ǡ���OF��Y�Q �@w�#�&�	fX� l��r��@!����5�<�p�8^ۆ�,���au���Ѝ�����@����J}F���n�^BD�p�vwvs5hU��.�oY�Ȭ���V�f�x�d<�9hP���i=�Bc�X�G��vL?�s�����u�	���p�TZ�#z�5�.�L��][?��L[���!�����޷���!�*U�d����<�q��J>��!ʓg�Ro�u�n�v�x���>0am)�X�o�<Q<�
1Үb�����+���*x�ͰX1U1�M�l��T��s�v���r��_!��G����eч�Em��O�1T����j}���P��`��]�*c�ÓeqЬ��Z�� �oe�lkv�Y����ReO���߁.�l��6�ܛ#\�aNI�Ç8yPx,�*U�a_��k*�7���p&�z߳l���j�t�
�$���s�7�Z��z��q&�H߉��	�R�sǀ#�����c�i/p(�,8Mu��Z�"�ƀ;D����|%�� \���rK��������)�[J��\P��ލH<��,.e��1n{=�P)%��Y �cRNއ�I ��<��XlxVHYEB    fa00    2c50�m�E�ͪ�O'E�y��:���m�l������_6#'rg�H��߽fh1*k��F��>�̔T�̗�?̜�1�F�MD`A�б�r�d��gj5�j bo�!����=+���8S/LaYs���K�U�Y���#�D+8�_uF�U�KE��"���	1OE�� ���E�_���is�3Z���~�D��2l�����r�s|�����p�A�b㊔�;�tF�z�����jƿ��
ڕ�[8�����fIg��̧�W�ݭ��S������� �4�"kK������r	����E���r�(�¹S���7�����N�YX��X|�@��_xQj���
��� io��3 �c�x���N�}��I�b�Z�m��`�h�>K%��?��s�-H�p�"��r*�^ۨY��|y?�?��@�Q�G%�!�(�F���Kx�*�˰�V_M�
u��Sq>%�G�O�����9���(jR�����GR���9EH'�<N�Qw"��@� ������뽃TB����u��@��'�ٷ�Kj4&慪A�$/�����P*��N{aS�N��`�����h7O!�3P_H�K0���PO��&f��rX���4o'�!�� ��X����5;au>���>�����H?�W�:���hCsi�۠�5hKn�	�u1���e�a_�xxx^� �v��j��OsIGfͻ��')�c�6�;y{Qd����E8�^���n�&�{ȃC4dз :5��7N�yH�G�}���'�c>��(HOVif]sXJW��_�(��_�(3�4�"3H䉍�!�����m�w~-a%�(��PNPQ哈0d�c�������(^Y����cW�f�G0CE�#�b��*�Љ�!`p	LW�Q�ܒ6�#�/|����ĉ��}^qs]Ҍifȍ�[��3Ϝ�����
>uG��~�-�N�Ș�����¾�T��쑐��kOᦊ���zS�j;��&:��w�z�.0<�Z)<�����?Q�j��֊&=l�U	��1��%e�.҄��G�)�.��-0�ӝ�-�sE1}`�P.��/�Y��0������=S��/��|[2TW��K!�Ȇa!uE�� 11"!��%+_C�I>'��i�w�� `���U��|$國f/�� �m;�#@����Z�^�d}��΄��l"߶ϘT7���#�D�
���K�;QJ�`@�Z��/�(��7w�CYֻk�Z�SbW�$3yO�-�[d׌��"^cٹ�CG�Md�Y���=�]5�ԟ��;�B�o�F�@��u��n0p�+��
��#m�'�ς��ۭ������V��2�PGLأ�ܜЂ��9�kǌ�k�&�7��v2I���������"sV�_T�1�S���5�3̶�ǣ��8�{�G���b�k;���Koy�b�,�S����٤U��^A�2���� ����I킏�����/�">�ʂa�ťw��fr+�</E��l������M� K�}ɡ9�d4�*T�[�dele6Q9����)Č�4��+���g��}_<���8B茺��I�tP<����u��L�Z0vy���I|G�e�d�B�=Ԑ^l"�b�O�e,�{�!�J+^:g˂����+���@>�I���7�0/H�e��Z�m��q�Y�%'/]�8�A.��5��nbQ�VI�A;?�%��|,���� �s�PMɈ���|��c9�� �������>K^b�ɜ�iaQљEî�"�������4�re�����}���o��������]c'��Z�i�����W|��mvQG�É���:���x��2VN��*��@n�H�n31�ڻJ]�F���`<�dMB���m��4�} �{]�ӡ༰��Dq�:R�Y�-��M�\�X����������M� 'mccS�i���r5ڐ�;u���UIꜾ_�N�����3�
Ѯ���A��+ 3�B�*�j��T�eX'ԧS��F��y���_�z+�vR�+�7{�@R|ck��UB���;"j�5t��B������8���^����v��W_��X.��x��U����u}^C����A�E;`�Ϭ����IDa`DkN��NO%I��>v�]/����Y�d;��@���1��w�Qw��}򎰖X�3���j����=�y�(�[��th�Ǧ�U�t�湦�E������Y ��/����R����,�cn��$��QJ��!���]4Jl}�i�ɂ��C�_���;��o ��/����Q�5��|��\��z/gC��ߣ�����F��ڟ�>��v86��;�ߋM:�H!��e�:5%a�U|��0d��z�' Om����|%{�">g��O���Fa����T"j�ka��7_�L<f����Q�C�ofnE�q�s�I�~^˞�סP�j]�J�&pb{`.s�Q�44�A 8kyYc��^tZ�Ka��M�s:�j�ε,�ڶ���]����]���ȟ�%�\VTq[�V�	��E��ڝ�����~;����r�����Fn?w&I��ٕn%��޹�~ͱ¸����Ʃ��aG���,_�+��#߲�"�� {9��p �i�����,.���a6��b'gS����c��(����ь0�e���<	cu>�@�<�w�P�����.L*���=�3����4hG��L�Q�rm�A���c�iJ�I�,3.��7V^z�����
M����2�0���'�Vp����KҮ��R�OF9!��2.�|�7g�����QP���8TԦXX���cH�B�н>����*,��. X�-}�B;y��؄��d���
��g[�p{�h�����V���f��QϿh�d$� �Xn#���ϥ���p[	H	;���E������k<'���n���1����B���̩H����E��Hp��)���5:�$�3~��J�N	�F�&�ZL�g1 ǡx �L�[��!�>8S���SA ��Է�[&ݕ���1[զdӊ�o�λ��ꂥ�����ر���)����]�;ґ#�����85��d�5S���A��GO�� �]�x��3�����Y��&������ن����$�3P��i�"�Gs��7�6�1{x����	�3��Ѿ;��,��q����׽ ��aRl;|e��Q���|,��l�������zj_d>� |3+\C/�G����Soi~FI��a�l|M�wKO��mh&s� ��Z!}8��`t���9N&�X������T)m���,&:��;�ߖ��N`p1���L(�o�UZ��\�DM�"�
%h��=�G}z!���?}l��=t|;`	�9�N)R��.��2��	��6�Y��Y �ǜfU�	z/��_� x���~g����tJɹ� /!I5��]p~'�	@�1�����T\��o#9��AV�A��1���=?2x�y��X�1 �/dPX�=�
��&3�������U�N7@�ۮ���FEg��<����u�{�TՏ*�����Ȳ/�ז�~!��d���r�#	��n�W�G�N��)�B��"�����읥Xht����JA�u�}Z1}�Ѐ�l�]|T��g8��1�?�lM����Cq�F���o+�\��_a��x%C�s�nq�~�B	��Ŏ�s��d`}oO���!�6ףּN5���/,ժ��%t����¹MB�>�������D m�fI��Oc�}gM����� �`(�Y-�|�@V�|�'�K�o�4~&�m����Wl�k���쏂��t���m�`���I^za��#�*{<lc]�#dc��f?@S"��	��B(vx��FuG�굤�d���ͫ��R�i�߰U]�M�I^;z�� ǋN/�=�0���[
�ӅނЌd��D��3�ً��-�t� �+O���P�;�>+�1J����F�~ǐ#�[�r�a�1��5�q����OH��S���!�_ݰ�OT5��"�Z����B/5"|/ĳ
6BO��(-O���g�K�1�3P���k��z��	x����!@~&�"���M=�����n"^!ȯ'���쀄�p@7�`��T�������ys��;V�M�`>{`�j�)�ZȢ��*� �F��dn�V�y��|H�����c���#��m��P�?��[:@]����#YI߹���l������[h�������,"����R�g�sPu&�}|8F�gS� 
���5R��X�@�`,�����exI<�]Å���''����)?`2+��Qa�%�K���1�z_^F#9�:IZ�ܻ�#p���9h���F�W����!�P*c$�"�D'�Y�3'��d" R��B"�ݾ�]S��dG�A~\6�ݚx|']�?�6ո�'~`u`�,)�[��(N���E���ka�۴V��l
����6�)�oSK��%hyG�+�˓#�ӯ3�����'�6�ɿ��͟[�������	�����(@D�Cpю�se�����]�{��jV�7�S~g�Jqӯ66^;��:&���XU&�"s�R�7̖Ր_��F��,@4>�
��e���m(�L�8�����I`�%��m4���o�"U����WΛ�U]��'�t ;���ƫ7�U��e�Ⱦ2�c��j�������<z��t=?���mvu�HtL��zcW)x�׋�.zі݋�6�,{��Ժ�C�4�ò�jj'`�U�Xh�� �p���'�cb�����v2��o����0T�$O:���c�gm;�57�.��7�Ő�N�S`d�W� ]�.������\t��!��d���
�H��%F�`�e�WJQ��Z�IsT�j�����;L݋l8�[�WkG-��_np��t�pce�P���k�"�s���O�M�((�(9�ɐ�[m����R�� g�T��Ϫm֔1Ow�	:�� sA�aA��X4��m�`4W&�� ���Ꭿ���l�-C5�?�h�]��
��2�<��23�1��J��h���bว2�-Ȕ��<�_%�����3H2�T�W���py6ק��oD
���)e�*BA�$����|1H^���Ph�8D�f$v�4D��pԳA�����6����^��;�!%�5����0ً��7�m�X֬��~_~奵п0�)��~��^��Ӂ^�y%R�O��1��#V�\��~���#c8=����b�0�+������D�C�a龎������^�	}�Au�Ʀ"k�pO���kKM�2/�|��]�_۩u�����]�h)��7q�tDv��ϵ6�FWC���R=L�s��k��9��[��`���	�*�0VR�,�Q�2l���&�1���J�0S��+����w�^��̂C��i�X�M�ײ ��Fӆ������]t�le�V���庿�l��w��p0�WnE���u�z�J�d�}ޟB�R����NKM��U��=°҇���6��O���_e՛�ms�!�eV#�A`'̞���t����jN�V��%�F��\�V��o��.i[]=  �jӁ�MIKOh8�K�X/��)��m���˲BY$3ߊ�n+-A�1���+��?'0dw�i{1E�}FQpʦ���	�U��%���ͷ+� �#��a�u����a2Cg�؎�*��1�r�C��?eP��bH�V���]Mo�2��v��?\�z�~J(�|��%�r�:����Eܿl����Բ}��$��ol�N��y����=9r6���)˰�#���O�4����<T�Ҁ��d�|��T�V�.j���{�]$:f|(Vq�����sQ̫�kv/�\kg�?��m&5��5ݜ7�#��1��V�i�ާn�z�0Ti��fVV��#�z�ЯM�����%1<�
����M�����K]Qۡ�Cws��Cp�x�{�Z��{Hk�x%��O�~aRV2%��W�j�#���l)��&썚\R�	/Ի.�޾Ae����A�M �m��5�nmr����T�6W�g��.�`�D
�d�1��7>k�ೡj��W$�m���
���|��k��o�4R�k�k��F~�E�]N(x�0	��iyY�y.ıNK!Ɵ�4��Z��>�����=)��­ط{/������ñO	/'Рnê�^�~5���q���4K1��yֈ#��Я��e;�<�}�zE�:_ӂq~�Z�����tԋ���͝�Z�5-,�p���͇*[���O�X��e��'B�S<�u�j��,N5��LnPL$�{�yԞ�Y��S��~��$|p���,ւ$��-�Y�&l��+5����qL�z��X�#�nWA�<Ԛ�u�*��_�%L�k�R�����y�����(��`��?�_��OMg��v��#ЬT�d��6E<s����t��[N�|R�{�_oW^'6X��׮�|n�]V��d�m2ͭHȠd	1�I�Icт	�	8������������v���X�c�[����`�|58����/�%@ƣ��p�A.�j8³CGCL���������u�3���_���Uw(v�G;���`����dg�h�V1�s�#��ѐ�G^ϾnZ�T
��+�i?!p�0��:�� F2�#z�~��̛2�s+�/>M�� �����[��DZS����ӟ,����N%1�������ᐻ�U�Q��Z\V���*�Ry"$�!�.p�t���F�j{~�)_�3c�Z�)0̿4%]b}��^����ˌOw�3�H����Y����J��vH���A;k�����<Heg��>��'���+X\��FJ�ȸ-��J��Z�蔝�Y��<��\G7��|Z*�'�<����Bľ�x��1�#r�_�уfk6�C��)�H���I���B8�ag6�G�~�q׶�c����� �}wy�k`�c��q	��2f���p,nȄ�z��J�����<��T*�Z[���^�d���|z��ϳ��{�̈́ Q�b&
�C�J�l���φ1_.w�&Q�ح�6�^�aÃ(��|,Q�&ƒ(�hnbZ��Q�+�!Jbí��S��֫�F�k?tzR#��FLU���+t��4�@`�o��9��ܘG�������}CZ�ڹz�T~�ѮC��)�-�M�Xq93�l���Ž���1jX���i0�#ڳ�p
���@WUN_�Ν!~0L}�_`�׎�T��g�*�ն5<'�<���_�'��S��꒤�)�4pqDZW��q5Sc��e�"�����[��"�\��4���ǉ�ԍ�<�@�A��IK,#�>6���A�K����6@�l�oDq�g�0��N�n6~N�8�V��)u��\8�)��zӾ�P��_w�'� ��d,�M;���SWr�V�"��r�?ٷ�3��-��~�dL�ȁq|َ�-<.�A�+(�PNQ-��N8�u�^3Z)Ɯ'H$`�P��d�}�PaD?�j�b�n4�|�y���	x1.Ҁ8�����6�$��:�A���Xu�^`�=1.d.�����@w��E�����C�HሿS�U��4��T�x	���I��tA�/U�J�%��=XW���8�`	�,m�k-q��.��`�q�`��������:�s�u6�{~���ʸ�&A��_G�0;,�j~Pʱ�� o$*>� #y����M���*�?9"<	�I�|�Z2`�.�X �(� ���)R�ؚ[XJ$Ϋ�;g��r�Ӱ�� .#�y��0����E\��mGld}���>M/�! �����Wĳo<t�?f��	�z�,��Ѷ���
1�f�#�|�Pr���O�')���K��s'[S���&��IjۂuB�?j3�/���:��bՈa{KW�@Ez�(�g�>�?]P�xI�����S̚�v<Ŏ���$H��n��ϷsF^�O��`E��$�EB	^��W�X�6� �+��xVJ�7!4���~�MtRh�]�m$�L���� �ے�o��S(m�}�$��[.3�xS/�j�W+*C@.d��pՍw<�q�tQ�J���ˇ6t;��v���%��hhR�!Drx�����9���ݸ�Pz@*$#��X([�L�wk�� q����nZ!�q9�{��()��\��|�����2ߥ����v*E#p{p�jظ����g�,��/��I����b���SA�G�b��Ў���yb�XB;^��m���()L��:��c9ڌ�9�������6.�=\�ݟ��u��r:�G\ya����4]ُ�I4M~.<��{aD�OJ4�p�◜\�7�Ѥ��z1GM\aI�t�#���Γm��9�i!��w]!| f��1|�д����F��y	�{̪�,����,���P��փN����=�[�^9Dz�����ʅAP�R��s�$m[1��	+��ot�c�(�d���a|�g��T;Ya��IL~��%��W'���1�+�H����2��	�I>�
$M*��#0�X�%�^�W]y۴D�����'k���H�qlwoV���:��4n�;�ض�w�lV]��sy�#�׻�]H���~��34L���済�!Ʃb����I����A�K(1H=ؼ�H̋Mr�Ȑ@R��Q�<(��83v�QZ��p���k����j�ås�2�NH�%eh1g�ԩd%c���t��ӥ�K~�#��^P��Y(�#k�K��\?Cr�I����G��6>~���.�jce����\2�@e�M��Ez����7l�1���jL����ϾGq٪\s3{YZ��]����Z��#��[�V�J a)C�n��e�$]f��A����k��HͰ$Rg�}���N��|?�@�N+�~�v���,��Ք?PMKʯ�R�1�<�ay�p�װ<q�}�2*�b9S�[��M"�r@�?�ې���gdү���V����J�U�Q境JW�g��_����%��\���ߝ����`�����ǚ����EK���cN�D��u�H��`�Paz�K����Z�8�
�V��A�q��{���DLѣ�.8+^6��"��\6�@��2aX��abw9\]�?�:+&||3�Y�M���2j�B�L��@k��d�hML����k��M�>��/VX����X
c�|��Y�h�nS9n�=�>��'���o3c�l����mCgH=�aqu鍷�P垥M��O�Qt�ˊ�C��2���xD0�L���E�sP~XJk���YA�BG<da�8cV��sk�:@�h�[L�9�.������F��/z�
�3uɄ27����y����
�	`���2���Yo�ao ?�z�\����<����3�����:"��G^���4,R�*��9D��vz�=�G�}ѨˆV^�X�g�x�s*h\6}P�.u�ж���F�����g�Owp����B��A�o; �z�p��/X�${�dlɔ~��H�����ڟ�<��q8���j, J�*��i߆�h�C@gd��;���꘡�j\�#n	�^�B���;Ďo&�#�@f��*ݻCd4�K̔��Y,D������ H#m�GKyR30�y��iq1�]�V��4����t��� ����Zб��4������o5�b�y��/�[Jv_��^��4��JE� �AIX	���̣��6ߒy!W@�ty��~6�Y�4�y[�r)s��u'J+���+���>�Dk� je�n�YC�!Ε�?|�T!�*�j�w�ǑX]���s/!H��>-= X�|ʍ�HL�1����.��K#�N?���S��ь&�TѩX��#\��o��%��Ħ�2�<5�X%�`m�U�=����E�������q.4���1�[gx�Eg_%k�#a7j�Z(C�x�nj/|�W��*&�g��έYxh{4���	wS~ld�O�J��A����Pꮷ��d]*�͙��d��)"3G�|}��_����>���/�����X������N}5"��(S��t���܂�1g���E��G����Xjny/64
���v�	�RxGy�1�A,�i
0�7�����ћ(�y�Ҫ Loyr2���;���$w=wHH�J�&f/H��yP	��� wC���t��m;+3�})0̹� ��5��z�πϵ���ތ[x�`��}��x���9sR�W����������P��И� "HpD�W)D���Su5�s8�����s���c�q�k¡����+G+�]�9��k�j'������huwʘ��<��VY�=�c���{B�E8$R�[���|�	���l>���/B�#v{��{H�+�+GIQR�4�0j:FQ'�<��&�4l�����E=���%(�'������0՞��x!��-�dx|���\�A��X�4;�Ҕ
��^���!T��Lt���i
���8ꅬt3H��[H���Oq�
k��'������^?4,Eʱ�ᵒi���]��}����B�zSu�km�V��5���%S�O�a3)O7�I�-4k˅����� ��{�zI�k��1ҽ~K�����M1�������o�lӲ|xl�q�k����-��]"�O.�+"�As~]���i�è����TmKl���R�RDp=�(x�Ѝd2aL����[��h����~�W��VAe�tb���\0R����N���C�u��޼ө�&���UAt��<�o샣J�J`@�/O=M����,�p�@�-���8�T��>�@����F����j�3�f>�!�r����lO�
*'��`�L7d��숾Q��V�OY���7�"{�N�Ɍ_�����z0��֓��3J�A��|J�F�@�,����|S�*��]H>Aq.��'���?�+l����B.W}��`L�L�t[��)����>-��Uԥ.)�,�0����6�h��U�t����1�;<��6"��S�����R.4������x���J� Y;��:�v�e�D@n�(�;�9�����U�3�Pǣ'��~�g��9��Uu1�:I;�H^��Kf���A�������ʮUa������� ٍK�^����Y/�M�N��֛��_-�*�F+{H*Б�8��_��%F�J��.�@4����&�f̴�S�d#7�k��\���ΦQmM���(�����L?�F�;�l��>�EB��1ݕB\Bl-��Nn�\)�r6X_��AZ�й_fi�w�tA�p6��h~��ݪh&ޅ��IT~'UXlxVHYEB    c397    2030��š���x�o�q0M��Og4��6A�����0F*Rk��k��"P���ո�O�����q��f����: �Y��tH���i*�Q���|6��8��ï�<��H<\Aw9��]0Y��W�vd+�e�=W@�u�[$S�?�� )��W�f���3	��#�����B�����\���d�����7���ءaN��n/�����XNe9�k�	d!&"헫v&ξ��7�FN���Tq_�*ȩ�)j F�1��5(u?'r��M��ѐs���1{a���x��(fb�n���$	��A�kVּ��&�JclQ��)�n҃b/�dt�5���q[�X1�46�s�`��������D�h���J�@��9p^�%�; P�X�� �X��v����i�Cqf︤9&i(d!fra��ԡaw�2���@7q�8ǫ«�A���
�څ���Ot1��wV'��l�c�g6�	��5?�b�|�r�F2pl�9��oZ '�'�C/��Q��������oY�����i;��S�aNV+�0@ �uQ��0D�b9���72��0e:�� �����۟`���^ܑ�R�����k���� ����dS���8��=� kx }�*��[H��c@�0	/E��,(,=ķ��\��~?��a"dWYvM�+�s[�B�ռ�r��$�������(��#�`_}G���0dj�R�w��"��]C��C���z����TV�t��/-�Zj�z��󩾓JP�l�μ=�����~ߵþ_,'�>?�H�LZ�"!��t���Ӟ#��4����FB�)��M"�3�c)��k�돢
�˪]��bWJRv[[ �s�B����_/�Q��%򸯯�_!����o�f���pjJ�|�����=�[��I�j�W&���pq�����f��::]&bt�^�b���b�Re1��V4�d�#�"��4O����C�$��n�5U���@�j�N��N3�e�V�U4�Ŵ�Z���Hp���Sen�[*=����%�Yte�b���b��f v��{焉������P@�j����)"
Cw.�6�y����.�>8�i��65�!�\d,0�ޑ3 �B�fp8�;�U_��6ȥ̫��+7��eVRt(�Vi&�;.# ���o���~	�q��U����e�J��'��m17������d�W��V��u��0�m�)�H��B�bc������)
�g�rC+���.&��BF���[�q�;�`���ȸ>&p�D�$=k��� �+?��  �gL�+��@V��D3
:�G]���+�H�*�%h+�_&q�����HaU��I2��%�Q	������Ou��G1��c�&��@�vr��~숝SM���2�^����7�!'�j�ܣ^�� �}m��45��2�(�A�`Ҵ:������(*����G
���-&z+�9
�=�eY��y�TQ񌶤�����3�*�X����}nǰ�P;��B"6��\�y�zc���lrBqٳ��A��ʙ Y�>�8��]*'f�����cF���oVh���!iWI��ƥ<xn3_���֫��=�4��C(�MS�Gя4���\et��ҳQU~���$���uCi�	
'9�ڼ���\��@����N���FU�\0��]���w��+�i������I��Ή{��<�6��ބ�.Jq�׶��X�F�s��o������t�F�0��I[���̌�(B��E ��]uJ1��y;�� �e%��+�H��Tb��G6¾q�5l��[���@lha�L��c����
]NM���K�G�79e�EWO���σ�M-S�;�}�( �ln�%���M17�]���C�
��0�Y�kI�#Sk�ث1h��#h�T�N�ld%�Lw\��h���k�����އ�Zk	�����g197�����%����z�L<��/� �k<��~�qo̶�>��>a����=���^R�߁����&9M��7<eX�Tl���ҡ?�j|���g<s쇩j#�_�6��\	:�\��c:a�>.��L^��D�����<»����{f��Yl�S���t�g�e����N}\�Y���M�}��Q�������e6 ��������g��ɯң�iW�+~ާrw8�O�=�G���4>���`���6�;[���A��*�ЦE�֮�;t9[R�kLq3��%�S���/:dhߑQZh��V}|��v4����q̄.�]�;�����/|-�@�{ȇU�G9 ���_|R�����+άN+�eR�����;Ry�hޢ����h�����dk�RG��sE!ƺ�Zv��;;F|��,�Q̽@/f8�D��B�h����zZ��Rm.�A�e?t[ ׻1�і��h�0��T�ԝ������⧲"Fo��KfJ�>5c��y� �n�(��Q��"?���.����&��o��z�b�2W�� ox!�6"�Z���&~ZsuC.3+�+znm��Q1�`���Af��+����?�l�b������֟�l��3�.kg���
΋�iF�s>��)�:m'�v=b��1�C�*i���"�ا�S�vu&K5�2��lj�j��5+�"��d,ߑz�{��GsA�#w�Ӑ�t��������~&�~o��X?�C ����ܪ8��?:`:H���a��N�w��>A�������k�#��7�SS�2�>�e���.��ut��'VǬO�`��
��a���(��P#�~zbY�N�O�+H�a�=�aj;4����i����!�=�,����E>\e�̬�$�����=*���9�a���j	ۜ�0�Ж>دN�2�]$�Y��
�;u��1�l;�?�2z��?�����R<��ȍ�l�99<h�Zx���� ����y5���W��#��HJBm80��OA��~��Q�6V*l�.�F"����"��;j8~�q	 �~'N8@'耓���՗x�I�),>цY��4��Gֳ��#���B�����Q{?��ުV��ћ���P�4�p��w������Z�_��3��̖[�X��S��"5�6��.��M�g���E�,*�n�R�_�%�A�2L��S=W*3���b�#tgSW���"�2 �b\�@�c	�s8i��Z7!��m��Q�����H�M�[d���">n�k�"4�;j탾�=a٩s_�]�d�w�Fp�Ar6\P�U�d�L�2U�j�^��&U��%=,��p�����*6��<~K���O��k��=p�/�g�s������n�M�� K%0}d�رy��*�6FgN	t'��	����CX�yx��zWK�B�S0.%�Y�/M�*���zvM��r��K��#��'����'����T��� ��8������4��.�#G�[WQ����{�������œ��^V��~"BH�&`1����%M�Ը�F͜����g��{CH�j4�����g
��;�⩸d3ߞ p�3�=9��߶�ژ�rg4�L�,�ܙ&߲4�9�8�L�jL���M�6cG����6�^Y�G��e�i��S���1oAAI�Bc�?�.��������h��f���ʓ=�[dܬ+Jo=7�o��։��C��APN{�����w_����d��U^�5o͉p��Z�/| L�����[�&��*e�Q���=��v��=�e6�f}����^ҝ��&����|s��a*@�Z��U�s��nE��Ɲi�r$���e
���g���_��� Hd�"��������q�" �c|���W�Xu6 ���7�v� �#g���LD��Z�{�,O]�(FvG~����y�$��b��HN$JR�t4sDVA�T��b��=K�����g��=� �w�|>�ͥ :8�&��xXk�&e��B�_����E�J�>_�!����k��~Ʊ�)���A�������p� q �+��>-4H�F؅�>W��]i�3S�O�PR��>�-��քW�yݤ`���+-�?W�.����GR �8ڕe��i��A�͒/@h�D���ŵ"b�㦏�=7�_��(��L��%�%\��6�ߒk�y��"ylb<�,;�+��t(ֵ��p����n��g����#0d�o�hB�ȅ���O 8���O���2^I,�Nt&��lz��D����mE�7X=	7�a7�ceB�6��I���n�]�X�.�����b�V��u���Pҵ�.֛���<�(�!Fh"��!�/|��]�y�F��m��|/4T����Y�sj��lr���� ��A�������  �!��;�e�6!��y��Y.�tŢr/��E��n�1���f+lx��m_�%���9t���P��G�^�s�ӊ9&I��-/��}�3��?��q�t�]:���E��%���$����%M�&c����]��I$���oӦ�������_ӶFD)���vy�Ye
�7�>��p�F"3�##��y���S����T�� �L@�4#��n��̂��H\�%�}�|��K`O���c� W����W�*���Q�H�(��Éu�e�����k�i��`l�(�p>�y�r�������>�_ O�GzCQ�kئ^���1?u�i�j�5K 2��mWg~N���nwط��N�7�T~_����P���~"{��8��V%��d]�7�A;3v[c�A���+�{b����������3{���C�MR'�>��p���m�4��#ɘ�`L��_㴯{��O���u��\.j�`j�4?�d}��š׿�	]U/��'9�9���]\��Xop�0���a~�=�g���<��g��_�{B�ԭ9{e�m����6еќ��&�E�.V
�s[�`UC~,�Qi5��t�a��ag����KM)A���n0o���ǵ��#��s��gU�!	��F�9�& mIb��-�ݐ���j�>�WK�a�C���rH��.R�#��B�|s�p�|�$菍?��3�B�V��N�%\G��f�S/��5T�����S�2[����oz�B�1���&����Kd<������t�"��s����P�Rf�(5�u�	��/��c��U�j�dNM�o	I�FP �5	�i֌,r$^�~X^�Z�����cr����2��?�ɸS�%m�_�E:��Q�U�m�\Ål�7���bh�B�t]�]ſ�f���~�h�yR�V���h����[j���w�~RB�>
/�BP����A	��؁0�L�g���M�
H��M �\�;��,=\Q?'T�Q7Oˇ���a�t�S�}ϣ�����4�?�A�bzX�b�oq�l�%6͂}H��~�E�u���z=�;8��X�*%Q0�b�����Ф�բl�~����8���PRO2sN�[��؂r���p�{}�ubv��ƶ�J��*B텟�e���h�Q���$����n��0��5'-���,[�����V͠J�JЊ�m�t�z�WE����h��0�L��r�v��R\�J�8�zi�5�I�k�}*B\L����������a:(�b�7� +7Ta���e�N�7J@��E�~�{p`܌�rB�n�e ;E�k�Jm5��=FU��t��5���Nzԯu�1���i�8��e�ޝ�O��F�a�ɀ�"�N��֥Pzjm!sX\�QW#�o<����9����V7Fn�z}#�^��![~Y�²�Jz�i�:Zw��ֱ-�����L����1��ȹm�1�@���P���Y�'����Wr�p����3Ժ"~X� ��zT���县Z󪰨(�At�����u�Z�1�Զjɼ.���L��*�:��5��?�`��ڧ��_�g��%"2�;����7hVRq�Ao�C*�jZ����j27j_!�@�n�؊�=^q����� �ϼ�ӪapM���!���_���{�!v���ð|�#HY�O�ҍ�ei<����L�6���xC�0-����8I��ǜ~�wp�+��]��KE� v����@H��Z]�9�IU�eJ{�;>V&ٷŎt�y���� o�!�)��|!k�ݏ�7|���Ύ��<���=Nب#	�N���y�"0j_H��ܸ�Lg�%-�!�ҐH�|T�}����>������?>9VhM!!zr�J���C�{��6{��/���]�`g�K����
�,_�R�N˚j�/U�1=�U?/i( ���ó�>��B�����Oܔr��C�Ю��拸����ir�m�,�$��	ma�+;����&��� �Iu�G>m!h��`Q����h4*��19^��Z����[x��`��?G�I���2�ªۏEp��5�[��7���+�E\X.���,���_�lVE�qjۅ��$':�wSB���=��͛�uM!U�#wK�H��j�kY����M�}�1�	�;�p��3��D�m��ǲ�%p��Y�aJ����h��^
��A�Z�\�
?�A�[� +�޹Y���Ql�� ;��ǦY^H�MA4]c(�[h/j���m@bQ�y<.V��r�V�;��&	���%���мh#&������Sx�LJp�������힦Ja�)nhQV��1��9E]���6��%:7��a��ZFS�V,kD��.%$uȫ:) �fi�ddE�n�D����P	;Ig�QN�1%��L)���Nk������b9� ���bBn��Y:�^�����'��d%�(�#��~�-v6��O�/���0��k:����z�e�rO�HԨ���s�����z���}A��\Ȥ�A��2���v�d1�x/�1��MX�
�}1I�D���5�vv=� WƖ���+ͷ���*�`a�k����wȏ�ȗt���z�+/1�aq�I[�ݥZ��28�N5���ط���X�$�ϯBy�Ja��C¬)D#�=��C�Uxǔw����>oo�<��I�{�Zߑ)J�/t,�z�bЈ��(#0<|�(K�d���n0|�-B����m	���Ī�졣�Q��w���r�jg��P+AW��ϓX��U�k��������b���ރ���'�ƀ����rY�+���ؕK�Ӑ���*&a"v��0E��ڋ4�
���](!�� gO)�fX{,W�4v���§���6���N!e��Z�ʰ�C�'�E�������G��bp�|y/�W5�I�VE_�I��J�<�2�3^o���t;Tς۟ct/�&jQ�Q@=���f)f�D�9�`��q$^�T1��6uZb61e5��S�/�˜e�&#`GnY��)��&Y�c,Y���;�҉[Ȭ��Q�R�=V�XG�s���b����eOR���,�a%�*Fm>��!�<�E�Ky?��Z>�W�7��ء����Q
ac�+���4�����:˸oK�([^.N��!�����I^�����7$K�*{^���{�� `���<i��t౰�"[k��[��=ܩqO�3���C��������<�` ����|8�,��
�Q��ڵ��r�1�8rz����� ��E2R�b�Ie��䣎��X ��A��;�YK<�#�J��B˩HA��9�d�_:~���X}���b��^%FH��� m�����$�����^�'�6hg��5ZNs�|�6��!�uc��xėc�A"Pd/��"&��t8��|qe�K��;;� ��]����(�M�8f��R!��i��Q�����B�@q����4��RX�rי}���|�� � �Q:-�`Fp��jt��i�M�.����Ty���y��E���]�@��2�'�:��L���	�y!?�8���wH)��^��cT�U�h��|��K�p�h9@h�*����(����i�Nޫ�Af�x4��]���^�3�=��tQ�@�s?�a>����lE<,G%�P����[� ;��u��<�y���G��4�TA��>�-��U�����R_Wtݽ����MnC��7#�[�G~��ou�$�����v+�dI1!ӡ��������0ɓ <����&���F�\��:�-��0�C�:v����&4|�o�����O+ �2�X!�x������M�����`n��4�����t���'>l���!�������4G�T��\�!�������<V�	T9�VVҒ{;̗�