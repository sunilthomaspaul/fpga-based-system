XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��H��i�\�v�W�;7�v�?����m2h�w,8����?=%&��p��/ϛ,� NYT�.6��F׬Kad�}��!`0�P��F՗�vնq�
�5R@�̝k��F�S7�Z�
f��4)CC�8��j����.+�g�Io�n}�~�b��y�2Xx���w���v+�:���
�x]���D��ӗc��F���읆>1����ـ��t��ꊺ�w��(:��խ�"���IY�
�z�aR�;g��5��t���@�ƺD�T&~j.l^w�xm�F/>�(��I��op���w%J緄�l�o��/�q�I~1o�H�tn�HP�w���4sK�g��g���(VL����h�pqu�)')]�8�7�s��{M����#V4ye({���[K(���	��"����e?lB�әX���u�b��al�}��os) �a���С��Dg4@ts3L��`�nQr������(i�4>�{�-n ,�q�}�����o��������N�؊�1��d���<�4[�����t����~S��cl��D�<�SF��P#����P�B)���U�,4)-`<G�}��;PI�]�t���g���	i����`��JF��F豻�0&��K��n	����]�j&g���A�j�ԟ��΋Tc�ўP�u�|a�L��Ӿڌ��
���C���)����B\l�6��ze�e�Хu;�( m̬��(���01����}!>�N"�� X�:��sb����y���"�XlxVHYEB    7a7e    1af0D��G#@���Y��[`�
i��1�!���Y���7_������E�@"�g� ��^�k43p,E�6�8�^M4��"�u��2ޞK&y�S��8+�u���xQ_#-)�]
�.�+^<��]i�W�sI<���z!xajPh)7��r~��2��	F]'�z����@he�C^�_1�~LFG$��|��
m�x�oM�i��gpo୺�>8�2C-AI3)6O��(��S^:��5���(PD��:,5s͟YP-�S)�H2.��3p[� ��n�`�f���<���MY��i��@f�n�B��L�&Qp/�65�Sd�T#X`���p}��ڛ�3�<��J����U����g�6�e��2���ː�-%$γ}J].(_&/�(�i�?z�f*H�>qB����ǲ�$9�ɮ �|���_!�x��܊#G�?a�S�������WpTL��USy*�r�ddгlxviW�,�x���) ��/�2X�(5�?(�_�R�;VW���]�xL���ǖ�-��i/8�V=k! �7ӆ��[\��`�{�Nv��_��s�f�q���j�-h~"�Y�#SH��O���R�LR^�̠��ev�~eȜS��)�w`�N�����E�8,b'�APe�����k��~�"����oW�ᣨ$a�\�>3�RKt������"�m�m_,�Y��G�&ٹA8�^m���t6Lb/,{o�7z���E,'i�ɍ�ڧԕ�WE!��-��<�����uv��P�2WRe"�n8��y��Bf&�F�*io���B�����-�¨!&��U��Y��53(U߱�q��&S�,5eF��~����q�4��֛�ٰP�Ŷ�\wL�?�;�<�0�ַ��vX�)���]��_~I9��L���ߨ�X�_���d�����H�O���E���e�`/^�5wP�7W�L��g�����Z�r�Vq/�fG�G���ՙ�a���.��h�7�n�C���'5��7��XN^��Ε���Z��$��Y2����-�|`v�Љ6��`�G�8B���]�e���p�7L�����������]Չ�.��٪␛�x����<��o�������L�c�ԁΈəp���������x!�e���B
 9ְ�#x~�����XJ�@>%�}=uۏ���hc�"��$y�;�$��<��ͅa�Ե5����A�I|�S]�,?5���sx�p6����5��g���$e�P"۸3,]��9 r�RA���$^�7��z4=F����P����K=��a��:l�;��YV�!m�Z��/-gб9]�P�2�R־Ě��!]y�oئ&�1�dYo�_Ȓ�zI�gqs��S�z����T�l�15>�_�bnnɺ�b��d��H��Sq�ʿ\qc�HE��_��2h�<ߴ���6a9L�����U�}���!VFF�-\O#�o ���x����������.��^~�#f]��b�����_���E��Jw4mÇcNTC|C����v�Qï�j"��tv��C!�W����>�Շ&�7���[tk��"n�yB���ZsY`�o�^�)��3������L)&E,{x��z|��>�[�徻�m#��<��U�T�)s$d�'�M(�@눩�M�1�+�8}�jx���li�}{���³���װ����/͘�\��s#"P��
P��!f)M.�����5�VŌ�\KW����������q���b��7|�n�q�R
��U�YK�G�2�+���\�Ӏ��=����`2'lW�(���[:��(	��N����(F�� 8�Y$sgG�&�N��n7��_Y�v�O_8|�~Ҧ<����@_�(:O�i�Ǒ"	{� #X.���U�	x�1�%w���e��A��N�b����Xް����.ڮ�=NEݝ(���Q�Q�[l�D���. j5 %@}��@;	�v@דq��W+fHF$�iÂM�/3o(�OS	8��B����3�"4���������Zq��6SX�3�0oU�u<���^�$��	�;✒oU�L������V�[<�$��	#��[
B�VS��jK��Z�&L1���s��`[ӈs�� �x4zJ�\�p_-]��ʏ��;��覝z�ˋx��XK�ah�:N|g�� ���u	���
�RC(TA�u�(�O>׌&&���Vs�f��QT��Ѥ�����O���Ч���}�W?~9Լ�?W�V��E��ivm
�ätcr`��t�/�@�a=u�o��[� e������3$�����ou�����M2���Z�q�|���Y�@�:��ɋ$�R�t�A��mC�Q+�n�&�d�#G#Y�27�fJV�O�?��ns���!~$��Ҍ� ��^����k0�3�8U��$����k9���Q�-�5�����A��q��0�I�qД�C'm���*N���f��z��'���*���i1B�Ɣ�v�y����w���q��z;��p��GK�0���>	�
;+p8��a�z��7�y����0Bј-͚�Q`�ol�TB^�Sϳɨ�OP�t�P�^l��̃)(k�����ǋp�Q{��d����u��lE�D��oū�	�T����<S�P�Doޔ��}��jw�M��9��Z���-��z���j[tP�/z
�n[9tmrؕ  L��_?/SF���h���w�j���[��"�j���e�"�)�J��eP���$~
��� ��v�)Ez� �H⶗؈�2m5hO"˖S24��{���-�μ��hW�Vy(=1�����q?�(��\�{%� O�,���d�2rq��\����L�� h�����z��ą�MW�z7Q�(�iD���<<��,�i`&�����t0z7�Z~��A��RA�YaL�R5 f�r n���7�#��l)j�3�TP�1�k�lh�ob��JϜ��.��`4�}�&����*ʀ(o��!�_(;F�c��E5;a=��a^�Mo>&�:�\�\MRV$�Vm��oS9��L��K�B���	�g�%���}2��Ř�w��濽P��eZW-R�7��
���>cn5�鞀�Tߨ1?P#��
Pѿ����l�4`�D´B_Iʖ�C�3K<8K��PJ�+��6ĴN/m��;�b�m� ��:4�{h��u<�Մ��(E�\�D�qo"5B�ܧ<L�g$b�⤥TIF
yV��B��5]�Ș�l�&��P��/�X�m}1Έ��S��of�fṒ�`F(e
B�:r~��4��m.S_�K3.����y�<6G�s�~=��Y��wa�T��?6�����Fx���34��摺��)�a���R|z������BǪ����
���)8.ސ�;�ȟE���eb�`s#Sw���a �tL���Ц��	���s�!���1����z[-�l_��۰�t'&���~QZc�	k�;0�k�=oT$ԏ���z��%o���Q�_8�'1s�86P<#��<6ϔ b�j�ARp�b${r����Zb��~�ܾ���l
�ue9�����F�Tsɑ��Ӗ�h�bǐ�N�ه!y�;(b2�K�!�I�Wo��Ck�+ ��m���g�u��6�:�<�ˋ�˦��+2n�����������*0o�`f_Q����^����X���o`-�qK��~���"�j�N�] N�<�*���ª0f׸^��2Tga�'\D.�\�o	5OfĎ�)�v���<լ����<Գ��@ybz����gn@魓�1���RgM�)��$$�)ie6���N�76���S���s�-��`c<;Qas�����:�B�0�EI�����y��ҍt脾���7��=N��Y��i��!�K����s\0o`��M��؝��w�4��0��ձ2 2���!�+�VO�>�/7��8J��[�ָ;�^ch=���g�!$� #}�d�����RB��Ԏ�1{���X�E�׶�J	���'z~��cv�DۀCa�%^4؝�+m��]�V��y|�6�Xy"J7�P�:<`��g��a�W�'Y{-�0�ƪ��g��y#$�`{��"���sl�`/��Hn�=Ղ���(>ߌ�F��ʲ��Y����9}p�H?!���/i}��ư��J����Ek��bl?�l��@H۰��찤���2uR��P�L�������6�X�ŞxǷ��lJ߮����,d+G�k]n*B��㭣YO�2>Z=��Y���3�������UMa���Ġ#���!]��2�ђ^���RFN�Is@Wa(m��3l+*���>��9���t٠���!&]��<�L$���C%M�Tlw�T;��{��7o��p�N\Gx,=��L�g�sy�;^�Y�oTG�#Y	��^(��z$�i���F�;rwr��g����ȍ�u�z��}��Du7�?��o�,GF�9`��~�d���>$:����D�N�0WHhC����Kz��Ev��,�Ϳ~ix��2�� �Q��2�r���_ �F��U��LT ���1���RC��U�>a��r^x'Ti�2Bڀ���t�x�+C.�+�`/��E>�icߓ��Ɲ����f�6�he���c�F�y���+Ih{�D�tb�ۗР�$�rtE�@Yӹ�>_'�m��ks8���c��	�B��hH�	���s��C?Du9c���z��],G���i�=(W���@�Y���|n줻�G귛:O	��d4�����*���ؼ��#pR�J'�Y�C�㽈��h?�jj��4am�΂�m��I��X �UT[���D�3��z��c< `dL?`�����6�A#�B�>��"m�.�j`@N�k^�}�Iϗ�WX.�w��FL�ZA�Ug�X����v,�O�v!�Y�봭�
ڣ�Ѽc\�O3���:����W�D�+�A���1>f�|�}�Z�}�V���-�y��ÉWn� �A����k@| ��W3���L���{p�����f�a|"��J0�s�ڤ�{}4E�M8|>��]+��r�2��̒�~���B�'���2�����v����'l�Z�E�%��g]�l���0=G��ƾ]WzrPј`���e{��/䒺�~�1U#頚���dù)�-�*�������o�[��^@n��FcxF_C�$i�n #�H�gg9D{ [� 0_��K;գ��Z��	_X�䌑��$(T��2���MJ���u	��=-�a�����|�ܪ�q%@sϔ�>]�#Z\��ڗ���ÉS���F�1�%fjJv	��6�Z����W�I������Y@��vƉ�
v9�XId���s)J�LD�U��sk>�Y���q$�q������ k�A����6\�6��	�$�⫀���xY�M_��Ը�_�`!�	!�*m��U��̓�P��残g�waK3�`gI�^�"�I�d��6E7Xۮ0C�+��%i�5�����_��1b�5I����5��to�,.R�z��f&�ߟ5X��X�@s�^������ĝI��S!͢�|�J���q1�Y���MP�ͼo������+��
�" ��K�PƏ�e�
��H�V�.$j�!yI�F:K�X[��Da�`ϳ��i�PDY-$��A�>_�2t~����H=�(��/�����AS�����o6�KM�qЌ����o�^��R����{l_�d�YR���9�S�6n����򦜁��CAX�Չ,3x`_�Mm��a����Ȫ#B*�0�F��M�X�{��1t�%߸؇�k��$��jf\��2k?(*���qx��M�V���^.l~��B|�jY[��]v7B��=��z�VBA���d1%K����r�[5�roɲ�M����
�T:�?u�I�w&��$-'�`)��q���p��e4S����`!�z�1}$��rԼ��0�,��W[�eR�B3����Z��~��������̢��7�֯J��pe]Z뺳�뀬���t�]���ʬ�.��_*63�qrGq6�=��o��Ś�����p�i�5��}��D��@Qޟ�����WN6-��;�ٝ��J`��-\*i��������q+��m�OZ�zT$�8�r��_�,�~@��ܗ&O��#�^��C��?�>U&�;�2���߳�0msx��ڌHT��y垠��� |y��\=��ܪ��umD����։KqB�ڔ�� �P����Mf�3�Q�_�a����������7�����y���ҲD7��R������W�A��ʻM��.];@/˾�����9�&�s�(��{-��	ՑYo�ͳ=�g�t1@B�����D���e<��^��I��"�-�@�Kڷ���aQF$�ĺ�2�E��(��^T?vm�_��N��/0X�54H3%hc�w�U�n���$�{�瀮ק�tIrw{_c��u��t
�@$r��x�:�ܖ�8��CF9��}.�D��?����f>�I����m���g������ T�����&W��/�F�Aɰ��
��33��"F��^ꄸ�(:2���4"�����U#�p��2�bSB��"z��^Ğ��[g&�\��o�g�V�B[R�Ƶ{�'2�x�e�ҋ"L�>zl�A���Ky���j9�,�)T����Vb�l�NC�qTb�Ds�C��W�)3}�B�*_iYT>`G�7��!e��bF�{�Z�q���4�d�.�|q��W�H��s�I0>�-���K�#��1C���(�|Ayr�Z�����Rp��n^���
�r�$p0��uyW���hi�\��.T�5h�����rS-�U�-rI���
� ̀r�9_�΁Ė��