XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����%�q�QV ��=�6�C���4���q?�����t8����`�nh1����ʼ�����%��D�rn��MV�o�Uv$�Рë�Sp�pmPe�7@ߴ!e��s��ͥƱ�8,�˱mgߡj�u�}��`w��tZ�Jֆ�.�w�R'�n�˄�Gp/O�V�+.[�6�k����ed``FK��K�ʈ-�z�9TY�͞�n>�͒k8��-_~�ϡ>��=�a��>>�6�Q��ն���_ ����և� �#q�&��D�H�<:���P�L p	B^W#=v*E�M ��4���_a!̅�S~�1��ϒ�i�����pYI��mr��u���:�x���ްa�3<k �l �p߶�p�0�T�;�;��u�����A_���<�_�Ώ���F�t  ã�cf¢��z�=���s�΢W���,���'�Y����*D~;(@�~r�dHM�q�k��鍓�%G2���lE�'��'�Dn̖�n����IC��Lt��?�k�4�5�_hg˽���������έ:�6�NB�7\Ii]���Id�dw`�����Ms=��Ɖ	u�Z�D\m����`;�-GS�n�[�$^�h�I�u�^%�t�����۝�nԷ��I/�d!E��y�9|�y?�S��&���������Ǧ݅\����$4)�����r�ן1�L�s���-����V��	��vϸ��v۬8�F�4��6�1BL�~�W���.��[nF�MXlxVHYEB    5fd1    1710N���Un�@$��y����j�� �k�c`*�W<Rဿ��.��8�r�ټ�lg�^�F?kP����W
e��!-9,�z�C��U5�&̅��4@m+�9V�(�8z��,�1�������?�E������ƿ�~I�%Ȭ�K=�n(�>$�{���i�����6�����䘞ΊZ�0h,��Ĺ���������h�λ0<���dY�ܧ��#�
����)��ҭ[f�дea��tʯc��R�"���fK����v0�0S]w)�A�h��$�Ȫm�5��p�� '�wo���[4���)e�N�M"��
��Lڄ�t�l��?G���U4?%��A�OTl%��������%�_�'+&�V?"���ۂi(ҝY��"D�uz�6����BV�'߃f�z(7��N�jb�U6%����Iӛ@H�������(T8
J)� Lx/ ѱ(��u��{t�Y�!�5\�ɵ4-��1���<�M)@��/p�H��7Y��uT�M�с�!��t �I�e�e�,~���{ϐC�8���׽&��3Wm�[^��3�����t1�jޠ1��[Í��Fٷk$ZM��)�g?B���7�-P1�6�
��t��X겒[�;b�-Wu� �b��sU�����׹GŦ`�I�WhwSS����[�eO}�E���fh�E���s<7B��Z�R���9v˞����6����k��ܲ:$	*xr��HJ��5 ,[�X��M\��-�|A2��,D�U���>H��V,�7��ݭ8�D��d�T�ʻ�3�e�y\�E����$4&���â���GÁ�蕪����ؑ��|��XHb������o�ɫ� 8>V�_Rnp�(!�m������K�q�]@����ϵ.;�ySq���r�ǲi�ǳ�Z9,,�s��/��q����hs��;&t��)�ls�:@ג���"�����+�c�]���w櫙�ǋ�R܃u�_Լ��p���e5i�r�3H^6�f~�Vn���ek�H^�LQ��"D@��`�V
$K�#]��j�H���<����wpf@����߀򮽑���h�Q���F%�� %LTxtF�hC*�K�a!�F�m��l�dC��,��{�=(����c|���	�֡�S�S��3���	��QIܟ�U�qyJ�l7`N>1z��&a����],�U�(&�2�	$D<�n�9�w<s1u>P����V���Y2�����<�=��l2�\~n��X��ֻ��%R�)3h�-�$�RXe3�L��mʗ�E�SN����X,p�O�Q��_���1�CM��4-1�x�ى��7��6�����	Q��i�C&n��D��8-�tT�Ŏ�2�7l��x�p� #�
�����5�z�B�;��$�h���c��-;#uà���R�� ��-6S*w��'FGy0��*�!�s�?���rz���q���&��o6�)lg�����:m��M����o���j[<�F�`
?l������W ~bg�{���QF�zX|��������A��M�?�Ji*����ոl~�Wg�`.����6dp�8��ٜk�g,�Cϔ�G��q�W;و����ؑn���µ�C��e�0�����}1�
���Yd<+#
:z�WS}��l�~�;S���	���u���0BL?%e�#U�I�K�(�Shث��S�������5�(�q�w{_f�ӕ��\�=�\�!<;$b̮h�J �"u�� %Z�TѨ#bF��Vl��t���o�����Z���P�l�RW$�ҫƩx-:�3u��bB�;;QNzydkٷ���j����d\IѼ.�M�q�}	��e�!�
�ͭ^ ���t>�V�j�eb.�f[FYp-'VXUf[�C\��"��7��F�\&n��x@v6���M��ݼj�d�+B�u��}")���#r�g�}��~��
��"��95c�[��2�B�����$Pw�7fy�iq�����@���ﲒ�b�! �C�ǆ���;{s"�J��5���W5��e&��NU�.w���ԡ�Yr��99<O�(Ww"��%�_ӰIIy�����W�݃�8 *��WT�U\-5V�ٿ��Ñu� w]n���\�o�3�Ȍ�DuQ�|��8�n��b�-̵���VʞsD|KvV"��z�F�pm�Q)�SS�l�kJ�SpsL�0�nK�p`b��:�6q����4��:��{"z���=<�*��oys�঱"�s3�
�Ix��T�[9{�ǄsKcp�ޤ����FEjy��N/D-T��m�`"�H<�3�گ9�ɜ���҂��,U-��I���T����V������,f��~C�����
J��E4ɚ"�'n3�\�"�d��2�$�}B!}Bq(��F3��$"���0�Ť0ߺ��r���B��|
Ӧ�(�){��d��K�����xh��	k�		C_�T�cm!�ض�&���� NL���DI�H[h��O�����D�D�X
���1�H�m�d�@F�77������rŸ�Z���Y�I%Koޓ��RL�k+�����ez	���6) Sؓ�yM&�LLz~E������g��^��s���K����Cx���O,�j@�} ���tW����l�2�����Ɏr����|������,yS���WEH���˫2[B>9�?�\9mtz��H�IIU���*�r�|.�gN�����u(!$LQj�2�?y1rw�>W�O����K�z�(yD��5�.����DԪ��D�{Q.���r���TwYx,��\�6*F8m�Q�]ڒ���(F�@�����It/�Z�����%��v2���ؖns�<|��m�[[��Wbqt[.R&��$�&Hz��ӵ.�]R�")]^V�>�Bt���a|��<�XKgw�]�`ORU�;"�;����߶?\5䫔.;��<�e2L��0ۤ^�B`��2�٧'�x��H�yBK�ߙ(�~@ �D��j�8��d
r.a�Z�عV�#����>lZ�?_T&��NuH�(�ο�[U��T4������P�H��zR���������[�� l��&�{_��F�(-��2+�U<�+wj�����DD=�F��*�H[��ھ�9�}T�r�z Wk�#��(�*�
桕�1����[�`��D9p�$g�R�V�4'��2�����R�6�;ֲF���*~��g!��Z��Y�ڥ��F�x�1�F#!�8x�h�g_�����b.���|��XL�?��T�����<�]5���ƨ��m��CbόW��n��a��l�L�A��4s��V.��1/T=hmSSغ��&D�c�c-���x�-�����\��a�w��Z�`{
Z�haq�~A�:��ѯ_B�X �������P�χ,Pʦ^h�J'�bB��JW�*c��1p����2XX�Log�t���\p��|x뭞PsG>~�V��𷉀b�^A~�{8u��3�ϒ~�֕���t���++�؞�i^�����e1N���[I�)I&$��D�F>7pw����џ[Y3k��f��V��-]��:���G�9i��2��d���A�h����t�,�Z_4-K\���L��G�/`da�'�������A�`��cB;���6�Á?FFV�������vxA!�y���n]�u�R��_
��A��q-;+޵�8 q��ձ��TjQ��[I��e�:�l�w�z��Zg.Fߩw��.�;
.���������F���3}AP�}���� �>�xI����w��A�̢Zv!;�6�����w����C湦�:�axC_�ɵ�w�������o7��k�e2u0.(�X4z�~��e4��EHeb�%�N�Jx�21yT�#�JG|�&�d��Z԰��=��r)���.U��1�i��g7��W���*���%���b
�����/ܽ�_�XxU�=C��3�ϑDs�DQ�re>���	��	P%��T?�㊄#��q����<U\^��8�+}���r���#��<3�t��]H'@F� ��0��W6��8��|�8�A�{$�`��L㑇 ��P�_�^8+gB���xR�ֶ�׸�NF�P�J���U�
g� �U���1�=y7{ͭ渨��/��|=d����m#t�t!}3rmh�������a&�� ��s,f��Q����h�*��Z�L�cf�����x^�ANt�U��͈kp��m�j@��A'[�
8��Sr�K��'�`�_������NA�#��d9VY�p�2�~}R��&R��b���aggx���ek�z!����A�ɏ�h�T�b��i�t�16 �f�fWa"��d�����%>��&DP�������o2�6�e�J������bq7fHT����a��l�U*4:$K��@�50�և�#�^�1[�p�E��Q�"O��@��Vz��~Y����<�X�.�粯�:B~�p�i��u$�XkF�
\���0v)��K�L��l�L�aG�,q��Ǟ�vj-b��b$[/���,���PƖԄ�.��R��!©t5�O��o)�P�Pޞ"�YQ7�ȯ���1�,�ˬ����C�{�V��|3͊��7����b[�v`�8<`�A1��~�d�S��� ����k���2��U�� ſn��o֎o:DT�	�M}|�em��|��8\xAI2}�*VB_%�%�NM�Ka&�6��f��<����cr�쉇o�r||;� @�E��I��β0��i!M�Я���	�&���<�-��I9hkv-�!{��*�u)�d�s(V�r'F����t�ɏؘ��8ԫ�8���'�,�9_ K����=pث��fESd�EwU�YՌj�ޮHƊqw�����,�d!��������\O����ێ�X��@�	#�D�(���ŧ[&Ʉ� �ں�}I��/�/�e��d%�"2��f�Mf/SZ�h�i��@32���q�. �n��:x�V�rS[��>	c�q5�L�
�m� y��5�����2Z6�O�kE[�aD!���7����!!�Ǿ?C��0s	�8���5�����9""�x���ٝ�9[�&�~DP�����Z������:�^��҈g�$("h=\����'��Ä�vH�qa�yee����v*?5�mӥ����M�J�����ۉ��q�����T�ƾ�h�]�āU������I��/��2-���)s���?P{Z(�Qۅ�ld��[�� ��;�{J�7�=�wc�\�X�.�?�d�L�f��͚�z;i(G��N Y�U6�D�d����	�y6w���sѯ1^ٟG��߄��yG��R��%I��� ��Ҧ&G�3�UE��:Q�QK���v:�e���70�(�8���g��O�qw�k���XEn���r["��'�84�~�W��.�ǻƻ�N̴����md�"��t:VZ0:�#�2����S�Z��2ºwx���JwcvBZ@,zr�œHH��ݨI�5C@����@j�m�_�Z(V=�jr��.S��^�2QGV,+�K�G>c>@5�L?�!lRBL$���Uj�y��ߟ�O��ᦻ9z��?x�P��D��;��H^3J"0bVn7���ѭ����T���9T��ތ�Y*mĻ�A��i�(�t�#M�H��RM�K�si4�w�u��b��2�_�-����L�!��C\�2���/�hz0�^pR�}v��<�N��H���m���zӆ�����C$�=�0
p,��b��'�P�K�D�WE�Io�:��T�.s9��?ՉKv�D�r�]�Es>5�Vm8�e��v]1�3�T����"r������!�
�I
s*����%-���g�