XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Wv��ܺ����-:��ӭ���+�K��TS�~�=$��&%RO(�c�1N��������V-�[��ń��pG���;�{|����$�$��~�%p��.��<�:�}�8z��5��o�$�8�{��?�����j����*N-G��1��h��C�L�Q1���=�lԏqLlm%���c{5HQ�\��O$�X�!���K�>�R���&�W�3[*��r�h��?#�V��/M��Y^b1T��}wn�+eE�6o� ��1�q�S�4��1���� �.%2�s�5��FV��:��a�b3��iC�K����� �N���0m�LǊ�1����	�<��t<?�o��{�G�zYpgk����@���/ZB�`�=�۟J���X���� +�wsR�;sK�Ӏ:�s�ǈ�����hdO�V/g��`_���'H;	�9���i�t�^�&��-'O�WG�=P9��1����HaH�Qc!Wj�;�#K�[[^{ƪ�W~�,�l[�u���X������Z���Q�-�k�2��C�\�%ħ��է<5u�����;[�,�|x�5�>)�%��a�1S͘���p�X�W��f���+~P滝����H8kJ�E��}V�Ck��Pl�)�jT�:d����)ߟiK�4w��*��sN����yq*���^&-c��Z��h��B��$4�>] CB�$�����Tɐ0�ɚ�3��M5�m�99Z����
� 1�S��1���XlxVHYEB    2327     a90��B�^G��!y�K��ӭr�F���v��|��}7Q��cA�g]ˉ�훕�1$�E�q��w&}ѱI��ў�@�t���@��i�����]l��4�j�/�B�@�H���S�3�Ja �+����=�J�Z��c#��c m*�jM���2k�'�] ��y*֕2=(z�����h���CĬ�<�L�B�T��Ν?��B61�މׯ��P"�^p��`��V8�n�Y�f�מ��]ܶ�W]�����0�1�c�6$��c�q�p����Pg+]~�0��I𱂯��	���Y��jO�ANrQ��9���T����2CqռCYd���@j.���kX��29,|�)P��y�;5Cʮ�bo3=�2Zzk��\��<z�]	�!��U��r�=��P����|��4,�I�h#1s�@���!�7�l>J-YA�������O_tK�.�@�m!�>՝/��C�<�_�=h9���A@�zI/�˞i]�t�֋Eʂ�U��2&�8�_��j�$Н|��BM,�89G-շ��8���+J�t�Sd펮W]�n��0<u�0V�]�|l��m��J,[u�;68Z�v![���V5���9���7Y.�����& ��Hc����g��ANl��x�9;��Kaz�GTIS�'�U��	&Y�&sj1��˕O�ͺ`mͼX���:�t�A�����a���G�##i�\5iQ�XA�uGH8Q���`��)1
���q��)�
d�.���B������!��|�?V��Q�����`��$�:��.��j��O{B&��2E��^�]	�AO+qW�}��YD��������G�ƻA�	�Cи4D؇:�@Y��UjO����Ն�S��oʠ2H��քpU~~?� $����ҿq�oaRu��hh�FS�Ѩ ��'a��<�9i	1o�	;���@�yA�~~��;�����u�Z�*� �i����I=:�Q�@�Q�E��Q$x�Ƿ�������[l��n�.�ʄ��-[��hḃh��۟z;^���roC�^ �gw�&���X���U�Az8����,�ұK��Uv�T�1yP�ր�<�@�#D�	�o�V�q�F%۪(U�V��~���fo����fɦ(�Z�������=/�&웇��7�z���ٱ�����Wc{}l�#�[��s%I�/]j��c�M\Đ����PR0:?d������`���4F}��G�#�ϙ�U�Hw�4k/���!q����7�W��לl^�Џ����ա̱���{������Vh
���f�A3.a2��V��E�-q9��-z�����"���r��4�%0��4��ɞ��� ����3�[�B~2�|�q9�@�����4\���;~�Z�&����{[�n�μ�*���r�3m���D�,�}��Tqt�7�o卖�	LS@���"d���8�0� 
�E���b�<V�Ik�U(�
qp�G�@�[��{�+s�%>_���{X�f�6�h9j���X{1�,�/ '�t�\+�`uX2�;�*&,x6p1ɹ6�ɰſln! #���21�����8��ŭ�~'8]�!�N�*����qک>���֥r"x�w��2ճ �y�KN6P�33W�z1���a�����I9�:�8�{1*�7w���W��{�$���|Wg�2)�����*����� �!֌y'i��K�1+
����ϛ�F������&+�t"a��x>g��+E�����$GH��'vQm^⬵ZV}0���%gVc�tn�`����`E-I�bCEJ��T�G���DC_������n|e�2]5+N~�hy6ҟH�F�"3��ǫ"Ot�p_j�h�<د�W�u���f#l�_�֘%3���y��.t�d`��᥁����{(���
������D�hˋ���m� �E]�F�;p�@��(�o� �p Wu*#�晅�,���V�°W�$���� k�4s����ƥz�YcE�Uꋰ�ԁ�R>�����ոf�kY#mq�A�K�>w�h�١<�C�8]�ь�JV���;�Coo2�=4L��t��=�*�
��8��DJ6ك�Wd��$K:=8���%E���b�-�OFΠ������<u�C�v���#�>ثf�
��=�2�9�y7��I��L|E�N�
b|�2%��ѵMm٥a�,�i��^oq���錮1lH�ydHi��2�	YF��Nnj!WV[�A��~�F�z껀ˡ\�CӶ��!�}�.�*i�m��d�)�m�um�W�����{�7ZA�ݣ!❪�*uQ� ��H�MB���w��|����У�>@D1H�E��
�.�|ܒm�XW��s��P24�w ��t��테iDw�e���	�$��`���9�f������JDt [��*z n>5�z�-��b�~��*2�}�u�����B�=ӟ,-Fͣ���K��>�0�SQCVs��+Z0�]�%w�x�*���J0���Ľ�d�3*��&�<�l�'��%'��������(��Hȟ��絻�à6�*�Oh+O�`��O%��x�A�@��AO���$F9�l� k�և�f������Q\��=�Ų�b��N�c��_��W OUgvE���m�~��`�+�rL拞 OxO�V�Ksb�h�sG�ި�