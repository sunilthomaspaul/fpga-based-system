XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��{�X:A�1���H�;|����\²Xxxu%��� ��W�h�-X�ph��uL�#�	�5��Vk����QK�r �\��UZ�݄�7�m��1D��I8z�=M��"ٍӘ�{P�S�k�O-6�e�����eS՗y���#x�nt���֗�>��-�@�1� ����a�6�$^�%��}�[�F(eR1@X[��n�b+���3�4~��u���޵��W�j�c�5o�F�:�c]��k���58����������cU�Ds*�
FIS�oA��*�5.5�U��mDȦ1Dn=���P&��k�� �q5��4�R�������|�L��Dr]�y�V՞�'�����H5R̖�K�$�Q^���Հ1�&�=� z-�������(��ո�{�f�����W�2�A�s�i 8�ir�$`�#LiÀrH�=��"�������u����EK�8�sJ�[T;����=��C�d􈣫.W����dV�����J�Gt����p���
������ʪ�tH���,Լ]�����.���t�vDP��&u�nD����S��tV�_�h��Hk0�'k^G;����!^�����]��L�B�p����.�k�]*��v�<w��ff��@��o��A$���`���3j��A�G����Gr���9G!�a"���~ө�e���{_(!����J~��"��`1�]���xW��Rm;��XlxVHYEB    38a4     d00D<3=���?���9_ɱ�rǃF���f�^��ַ1�T�?2�W�ߥ����W��xچ_v�D��'��~�ꊴb��e�@d�����5�h���U%X�`^�X�\������ӻw4N�K1rS^Qx�srw�;�ȍa�!��w��v����x�v�|c&=޹.R�o��)�؜�&�Vuf���Q�T�'�ګ��Ԗ���C Tm��,����v"�L������t�{��J1.H�֢웤��ȷsz!ԝ��s�[h�/��'����Mc� D�����v�Q�3T6��X_�=�����֑��ST5G�wTs2�^l*��jI=��������Rjͨɑ���m�3Mq�
��������m������������R�:��/��V��KFU�~��"D�D3�b�:���WVH�YVdf�A�/D�N�Qq#z��'��n��բ�!QKULC��w���ٓ�7~3K�p�:K�8Mz�R�I'ݬq&u�w��;��DՉ�c++��)n�C��yJ:4]=�j���G�hݩ�~���a��J��X����4�zq��W��U@����\�=rPU��?�5qY�F����(���8lw���#w�.?=>�]8��j��m
����d�� W��,��B�7��zy���cҿ�#�\2���s�a]�����r}�?5�F�wV){��e��`,��j⵾(�@�-9#{�a�<�Ҕ��<j|�]�jJ�|>7�������k�x�6������}s� wH߼��.��I��{�>v�¾�G�U?��M��(M���j(0?�h��"��_��<�p��a�A3_�W����J �c�i^�K/�+�W`���N��N�3�Y
��:�g�s�rL�CS1��=��F�g��:��"�S��C�=��g������ș��Ld�c懿
Ϊ��M�!�����{��_|2�3�rwN�	�+�r��	y���i99�ni��<4�vß{��+��2��$a?�]�Lf����MT�en}����ȥ8F�Vڔ�@�LT6���,����i���W���:1�O����Y� C�m����z	C�����
����}Դ�8b�+Џ���ec���A�3x�bw.��/
�T��%���ˋ����@*�~/e����O�(~6��j�Ć�J��uҲ���ڗN���>#>�H��76���\4���U�ޱ0����E����]�	��:�T�G�����^���d^�Fr'b$�N3��sc�i�M�(�P�WL?F!�}:Q_��w�P��la��!�c*��^�eaw81�A�֒��]���q�&7��D�`�F��i���:����WfQ�#��_5qZL�v����(@%� w�Z�̮u�*��yř�`֠��.����|�
nm �E����d �I���N�>�תA�Ⱥ{'���e�<���ב�B^,
C�h���/hZ��؞�3��]Z�m+���L� ӌ�?�lH�c��6ѝn��6�:!��A.�������'7�bhD�->Eib�#i���"�h2�V�MiLD� ,/�����(�+2ĝ�d����!>$��S%^Ӹ��K�i�P�2��a�Y���vF��1���z��}��j]8���G�����&�^/42�
Ҳ�w�fE���^T��ω����B�f<�  C�E��
�(�P����<��$�b�;�N��L���	.�Hm壿Xb�]�g�[�my����l�'�e��
��܌X�PQ|d�W��>�Hׅ��?�#��2��5���cU�#�xȁga/F�����b�3k��˧���E���LѠ��ދ˄h9��A?ѓ���So��y�<h՛�8NN�[���j��+�~�.�7��p�?�;��0��(oݯʆB�N>>�L��kM��=���Ja�8��Z�O��ԡMi!��?l���F� �+K��FXt>_�Ku�a#���6����j�}m�f;��.�1h5c�ֺo�q�g�|)46(�+!�������d���c�X��l{v�����g�*/�4P=�����}��u������cD�x��2���Ԇ:.�"�si?��*lh�1��z�N�\�m�p��ʹ�õ�m]51�%��;��g�����g�j$�*)���;�Y^A,��2�ӈ�Mt&gkV��nŵ�`��e�"�y��)F�.jǞC�׸Ɗ5�(���\��I��˃�\�:"�U�V�= ���3F�����F��l����J��-C{t��t��0b9�s�c��S�tv����O�z~f�8�q&[��01��AY{�d�_%oc���
^���K��fn��G�	:��];��ZYA���l�d�V�^@T�b��:�lg��:�eLq+Yq�'��dmi,��N�W��<��9M��>��<,���`4�⏋;�F�4<��*�è�,�~Arȷ�k�Yi!���?�`U��t�t�b
�6��y��S���7�^��u.>���;`˓��V��i?��K��/��!�z/�>l��e٘����Ĥ�:�Xf���Y�T$`���P��@b�Yo~�ov:y��x�vC��fo3̡���9�g�=�k'e��1����?���6��~q�zX� �J�̫��6?�פ��:�bo���P���F�����d	�$8Iv�N�\�B$����Yl6�谌v��a}J�QD���\���!\��mW�[#�M�@5F;�$��u}ቚ9��DMNN&޳�N�yfu�@��o؋�|4<��vE,[S��A�8������N0��D��^�D�Y_���v�c��r�Е����B��<֦	��o�}����$	� Q��%Ƕ�߁��c�0Rw�(.U���l�����ov�]�8��@�~�\̬!,�[(�L��O�ʫ�VA��P�v��if{�+Di\���'E���r��L3���fb
`1/� ���Y�����䲅��1�����R�wM�XsKtđR�Iñ���*ΣQ݃i�a�i��:0�\+M��ʓ�#V��Ќt#.
f�vJ�W��o���{�й��o��/��.?e���T��q��%xV%��e-�:�y!��!�*�w3���p	t�f�p��$�k�m���,���C�J���&��[�? 4 ��~G�.�͉��
V4�x��n�V��!�?q�}h�T)E�B�w'�ƺ�+<,ӱ���):�'J���8���FTOL��V `h_��H����P<U_q-7i��/g�$wfODP@h�a��`*��������-