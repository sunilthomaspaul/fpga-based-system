XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��,V�_�� ڈ�ߠ��8�T�`x����X��O�K֕�@�1RE[�}�g���:3'1�(0�����I���3ݮS$��B���5g�:���.w>smW�P��NY�>Ջ���q������{��,�[4�D-���OXu~�Lͧ�0��\e*R�r��A�8C�T ��6^�u��O���z��Z��3���[�,��;��*3!?��Y�g�ϏzXd�1�l{�	r�h�۠-���_�A�wSJi�jPT��lٰ�)v0����֥�+��KNa�;R�[������7���t���j4�������E��^�I����)���Y/J��xvv�ԫ\�~4�fSx��.m~�:�ӱ7�۶��=�����?{�Z�Փ��k�L�����gMh�:;�����r�	[Q!�j,��o�Z��Z�E��fZ� 85�ܢG{�6(���E��*U�g�.$�ݍ����G����L|0x�?&o��b��~fg .���j�n��h�6�6�sK]-�.��!%<ڶ���e��p5+�(&�� ]�����eE�:�5O�~x�ղ(_�vk�v�U�H�^�gNsA�&�X��`@��m��תߠ�b��KE��d��R��tCl�^z����,������a�L�/_5{��l9q�s�v<��4,=��w�jL?�t%u9�)���p�͍]c���6B�&]m<�*����t����?���;dA�\����J�'H���k KYii&��|PZ�2k��㔁QdXlxVHYEB    1e12     920�k_l@C�y	�Z�92"�s�D^�E�8�ᆀ�4Y*P�Eh����);3E�鍵u��_����WLU�C*چ�o'���:D�Ԙ?q����M��
G�������T�񮑋/��>������
�Vo�r��i%Y�7���_OK*�=�l�a���q@0���f��8���gMám�	g��z?-쏜���JW��\�,���ݩ�RڼԖ " �:H6o�b��2�YuvQH,�@��?4ˉ�_������£3+|S�8_'�[k�tXnA� {�kU@��@8RcN�D�
�m���s�dE�Y��Q�7�� ��T���ⅽnN˷�ѰŁ�n8��s�	���EW������?[]����k���e��NdP�0�#aV�x�9X����| hS����n�]蓵j�be�u�������Ԡ�/8�ĩV�&Ҟ��)4�>s��!�L��Ā:N';B��w+��1Q������M��Kg3	Y��^x��)��hfF�%9��{{���� �aL�آy=�#��߽�}2��c\G������$�I��9�K�^��K�Az<��x��i��`{&�W�{ /&A�.YTo@�4$@�-��qT��&�ZY��/ݛ�����N��@<`2ƅ/�Y���?L�cQ��&~���
�[�m�Uj�ZC�x/vW���Oz.ԈJf�p�Хh'4�o��K�r�t.a�8E�ϻP�+r �r��O���f�l�@FO��4\��h%�H������'�2�9�w��P��i� �g�^ۅX𡫽u�ը7|4�7�H�}5[��t�¥p�Jq^�:֍0�9c�huN���2�O'�-9�ԗL�a�p3�ŤE��&��t�J�Q1}lp�'V0��o4�wX1D�~)$Y��#�)���3���4q���%���~�߂e�S�dsmY�鹍�o��Ey���a$����	<W��`��-�,���P�G���A�Ny*�a3<rYF�e~5n�36~���w�4	��K���j�%bW"�Y�4�/	�
�MZ'"�J�aKX��[���&�_��������D�fi�9N��*�(8��j����ހX;��9`��8W$��%Ӛ1C׾�r�U�"{��?�.����?p2�s��\��7� 6��h��ޣ�,oã�Qø�s��5��!�'���9�Ρ����#]C{�}�4X�b	��*!n#O�����8?��(�X`ږ. k�K�$]�(PMe�螁`
�b,�f�SY��P�%_��N]@���g��8�̵w��0l��r��V:�'5Y3�0�/�c���}k�&�'K��?���2�׶Đ�������]DW��m�5w~�DCK��3�ኼ8�C�_��q��kՑ� 
&��~&��_#�I�\�qȫ�P}Է��� i7�c�>� ��Eb퓃�lA�O���I�H�'+�T��C3��tԴ3�dIfS:���PϷ�u�1��5xa�D�O�1N9qH�g����+�,�v�ښ/z��9[nz;��6�%�j�6t�ϩ��������K��$��d��/{����֔�Y�R�w�GL�yB���I�Lib�;8̝���0�j)#/���9cP����9a����qj?�N`֪�g�Cɏ�]ɮIU?�<8�S#�y��P!��o&zL�I,���޷o2~�֙��g��#��\b\��&?+��Iq���Hh�U Aj�ˑ��$���8����_Z��<h�aW�~X�����87�2�����^�8����^3�/�O�I+b ���C�:&�������-}82�ʶW��{��ǚ�
C#���-h6�$�1�\�+c�j�P7u�V���y�aoK�
{s[؆�+&�T���j����^�S���^m�U��*Gl��ps4���U��������~���\�B����������\�L�T�9wŁ�0r(���m�CS���2�����2�E��1���䬭9�l^�Q�w�C���-9�����3~��&�<��g����s!��~v�:�+ZlF>��zT�ܶ�E��v)/���8+�0a�+��q��he�+�/�C�������:}���i��+;��a��Aק�ft��������D�������ÜW샵}C�\m+������^���5�9(Nq,��u����J�+H&W�6.U���u�c
V��/p}*����ޅ��)~�TB�	�Y�ا4Z��e���{Z�>�q��%n��62�cfD�yeD�+�����^�`{^�Y�����.S��Cg�%�mX����_��	G����]V�^贊�*/��o��Ă�Y���|��m�n]\	�]�����	@����#