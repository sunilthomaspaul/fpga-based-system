XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��G��!�\y[9�h�^�sΑ��q��4b1O&ȏ����S����R�6VT�r.=�bд�t�N؈W��$�p-G^O�����!m$�]��r�$��OV&�Q#�lՐ3�v���[�k71��?4�28Ξ�����t@we\U��B�K!N�����=��e����w��O,9�*C���B����@8��m���fP��Q7��7y[~��O���]�3`�+ ���/��x�/�� �{Z^�/�n]j�K�V��r�W�|���c����˾�]l�R�'J'ByLKI�օL�BYh)���e�A� ��iO��B��I�J��#��O�v��=�uԋ%t�0��.�i$�2�-|ڡfW?���T��m�
Ү�ѭ{¿�Ɏ��-�b�3���)K(R~&��	��`X`|���_�'(M��@zpL�����������������jɂ���P�k\�<�r��ϟ1Tz���ss�e�9�짗o�]s?9q8�[,��g�}Q��~Oc]�~0R29��=�5��F�a��XV)���O0���ظ��j�v(��kN��@O��������f��^�;��W�������W�=qPrC&��mBeu�%eQ*�n�۷	����	�"�a�3'v�oޚ�?yub���9�(���$Va���9-�yS���]��׽K�c�������!!
!���5�̴T�\k��j��K����꓉��]x�����UU#XlxVHYEB    d81f    26f0�iu�����>]O�(Í�-P�&q퉺���bJV��(��
���EA�O56�/�+�t�7&[@zH�Xe}yD���:�S�Q��,�YR+c`��E"�x���֔�������bYe����� ��߈Ӓ.}o���љ������D���8KN�"A�wLl:�*dX�c��b�^��c �ڹQ_Cy��5�����2�s+������V��XƣƐ� �����&|�z�a �O�m�]_U�%�f�죐��}��C���ƌ
6�����XY����2Y�1���-ء[`��a�>��]v����^N#9��	��gE�Pk��$x�q6���	t��v�DMMս��\�B����{��WGQ,�� ��/���lj��H�%n�	�̈���EW>d�}��Op�Vh�\F5+1�zM�y������d1�t�`~�n�e����
,����U8 {��uQ����<�&�l�{P/�;���0ߕ�Ҷ~ #�ן��{N5 �Q�6�9ͬ��3�I��Mc����m�>�%Lc\b+єo92W����fXk�O��.�����(�̒����Ӈr�B16���J ��!�b,o���Pz-u�þ�!� G�iV[�N���ȵ8��j�ᦖ�������f2E�qΙ��X~��h�.;�N�r*��u����
W��(�D���Y� /a!�E�]�C�v[�i�����٭�>2:g�����Iv!��X��ϕ^��Z��{h����{�f;����x*�{���IÛ���wB�#�;��)��m]�9�u�hZ�*�W����L������)bB����X{k�Rm�̌Hݧ��U��0��o�w�� b:��d�-�@�GģQ:W\i�sg�>L&E�k�2�P6z�!��m\���)���< ��*橇B�6�y�۴Z?�SѢ�*B���G�	��������}ߦx��z���z$f�*�2nJ�>�v6�x�M���t��g��	��^�JC,#&�)�%Gݢ��4�ۢ��%�׳`��]���^B
f�,��W����/�*[V8�/\ +<�Κ��m�TG;�g;�=ś�i�%�c�o"N}Jj��=�2t�"1"S
����$/~du�S��}��	�2�<�зH8N7�"k_?�D���Yu%�Љ�=N��ź�z\_�[fn�e�sGX���ȥ?F�<��L�ź�sK�N=qۆg���tD6>��H�SDa�e�@���OAև�,}{�	� �y��װ��]��<b5�GʾS���K��	ڮ��3Y�&�!7`�[���DYn#�b ����ܙLxx-!�Ҿ�	��k~���4*��~��)���� ވ���*�!�)@f�<�}��c���E*�Ni:���.��9P��r#����妖%��&��7eE�����\?@��7��m�[��DҠq�����?��$�R�)(>R��Y���P��G�O����0�=^]t��T��zQ��<�1$l��}:�vw'jA�u������ye�`��,�em���Ⱥ��ۭ��3xBW� �?�1�M9wG�����7��[��� �Н��	�gބx��������G����%�J�1�!��5�� �V�*�7�?:�OgKy��Q�ӄK��P'�
A�H�e��E�r�������N�pƮ~�u�]0�8�������s�el��^[��6��t�H�_Fx���P;�]���P�a�;��a��#��}0>P��*$��Ҩ�H���j��4�/��ԛV(�X/���qa�I�0�rnI3�Z�����\XCփ�`���mcѶ��?���$�J�����]܀L��2��k�h���ZƠʧ�������[E۸�6�5�j��#�`4�ʾM:�+��`=��N<Ao�\��{��Np+�"�;�KRZi��'�|�ZN�����e��ܥ[L��j�m�@j(��-ޔ8N��첎w��\��$��E~�k��j�G,[��k��T���V�YR�`}�w� ����G
�/.N�o�t�J�`�:�^���C�&^����k8�L��������,��N:�U�T�� �
������/�4-3�j�+�2��,�����=����W[J��'^j�/���sT(Ii�<�:����.����#;��>.�Uusn^308����m��!�.AL
� "�D4�)�g�� �x a�RO�%�z�M�;3mr�)���)�Q����\����$�Y�)�"��岟auL�4�KX�O��^pdo2<�����gX@��QQ�F��j@,��3��9:c��{3���u;} n��T�6�W)����_^V̸�L垕4|�&��oz+N��� U�H����qz�q�����,��%R���Y��p�-hq��S�ǜ���+�5"�9#�l�C���<��&k�-�8��$d{Y�
DA�]���_��7���4M|}�&�[7o8���2�I`��/F�ׂ�$ ���y�J�Ġ�#C�/6e��%٬���ۢ>�3����z�*�ڭ}�[|X�.n�,�Y=�[�v����E#J�7���'��{������8g6	�~!G�6ܝ��.V#�ھu+ji_�w�ۉ�t��s"l%�lu��kBE_��R���q;(�6�����ǽ�ˍim�IC�_�/�o8��1ׂ�Ra��֝0s���y�t�"�Fk"a����T�Ğ(��lI6h�;j*���Ό�o=��PT��L���5<w���m��gA���A�"�<�;̋�+���о�
�e(|!�>W#��!�Mc�,���)�bcku����)K\K��6Xv�h�	)c;#����Õ\@ �B�D�O,l�9�#���R�W�� 	ق � sX��E�l���272���N�"����F��y�z���]l��A�(�s�(�{��9�9Ik��#?jS" �k���[��)����A�p��qS:�=c
G��uږ5$Tٸ�Ҵ��!�����c�q�9����7�~��=R����t�]�]��ާ
�B������]ϊ��,����`���?���eU���2�ؼ@/y��t�%��ȷ3E�&�ZJ����!�w��Ɖ?���0(! zD
9��7�R��wsWa <����$s~�nl0`�d��kn���h��6uo�lu2��
�|�}Ԗv�zIa��	ƀ[w��	0�*ʆ���!���a��3� �m9�"Q����gI�/��|����6�ezh!�:j��_*BĻ>���=U�X� �� YEj��TW�޲Z��R�>��������H�^�Q���}~���%��FH���DlF�6���s�g3�T���B����o-�m�l��'X��z�/�o�m�)+&�yX�� ����������.5,�l2��i�HE����=�9����F��bJny^��y�g����sS��@�vF�7�dg2b�����4Wkpq)�1��26[}s�^*�^��H���#���w�׀\������GupBU�D�	�Xg�`GoҬ����ɥf���ı�sxR�ze�9�H��B1�n(�"bPM
xSv���-�-���NG��޴�@i�V ����ʼ#�9�ZՎAN�\ʊT����=�R�ϛ:/ΜQ�o4��RӨ5����$��\?є�������s;��y�:Km�ee��3�jbӰ��G}�}7���ƹ<�8��t��r�&Od_u�^����Z�������fl^�pB�Sh{`E�Ѱ~ahc<$���ws)X@5C��#��;][���0���i��Mər�����kC�]�Z ��YS/�M��Y��o�s�K>~���~P���ȣ/�60Y6=��L[k�4��ؚz+��Z���f�'����̜Z���'�hX�0j�Ӎ�ـ1�+���G|�1}�Qq�J�LVju��+�n��o�hp
���׍0�4�':���:�|[r3>�	�<��� cW'�~��l�8׉�k��I��&"��܃�q�Iu��G��Z���V������_#hq��U���^�k��^�
�xԻUI� 
o��6 ���qh,X 9���xԨ�"�%�>�	�+���%\Yz!>r����]!�&ԥ��j���?Oqs������jAQ�%ׅޠ�o���>�����5��'��z��3񋨅��C�9�+OAt�E���<�N`�Rͱ�%"�7=Ðavŵ��5��5	�W���]�	�c�*�NL���w/IXte�{��%L`u���x�f�;�uH�w�`B� �1`?�͈7[���q*�!���O��(��gz5�+���]L�{ʖcedix�?�t��#�ka�!/DY7���9V� p��#!\JA�ʸ �Nw��3Q�H�.�m³b@<e
&\LX�A�Ӳ!�hT�J�r�!�'���Ğ���)4�g���� ��y	M�|�+0�x��?5G�8���J���A���g�����
bP"&8}�a%q��x������bGxU}LW����:?����D��������_� 
0�(��T��������2�U��f5V�� ���顪zk����!�Ƨ�R	�$&p� u1��ާQ�L��q���p�����lk�4�������\��mdL"�x�N�j�J3#R��`�Z�3A��ց��Ż���ߒP_� Z�����W���O��Z:�e{SG���ü�a<Hg�4���r1�&�Ժ���;��X=	^��a;0'�̦�3(DH��[,����w~u2z�Dk�����3 _2���:��i�.����p����Ͼ�e� ��o����l����u/-EU`��E밿i�lՒs����>�p'�0eѣa�i�!�h�k���.$��bP�8巯�]�Pd��+Hz������E?@���K��ӟt ~�D�%��� n���Ե�tq=�כfV�B<5�?!���~��{�=e|L�Y�W�Ư����J#Hi��E���AzP���J�\u�`8�3�cv'�قu6�4:�T`X�U�/�F������Ut䃞�x���|�qm���:Ԝqb�p�u37:�M�o��~�Ä`�>՟�53�5w��"��
��Q���{��f=��L�g��;8�w#v�%v�wd%���/;DH� �n�� D�l;3����F�zɨ�\�-�}s�$��FM����i9;V:v�9�o"'�4D]���?�&���!4I�R<�g��B"�r����L`B�I��̮nu���>��],��ꭄ_�g˂�+�!AR�J5ρ݂�.��8ſ	c1?7�7�v���$Y�e������SƝ�-�l�b-AP)�����3���*�A���?��
I�B
�)�N���i�|p�	s�t��T�%!�h����Mj�5��	�bj+���"��%��Y� ���\��<�HYpU���K�@K�z7��!G/{تP�MRQ�B�cȉ�������ob��� �T��)�dgjR��Mlv7ZE�f)n+/�wǏe�ڰ���s^rKMJ�|-���T��@I���J�u���?��V{�:I-W�hn�%�l�#7��+��Con뀝OC��Z/�#�h��|���p��P�ƽ�����6�uӋ�<^�_���8�gc�N�ufo�F�|�=)���v��zxN&6?|�m��7�3K�c �qAM�p��7�+�U�%���)�]d.lj𔜐�Rͽ�r8��+`���I���xPa�\�䡕(�ꌈԮDNf�G15�4��U�0�,�uM}�����R����g����b�҆�v!D~�ebD�E�ӄ`ә%�:0@H)���8�H�k^&��m0!�j �&"�<â	�gpm�pz�[��X A'3�t�LXi3_�Ք�e�!��_��lĭ�*�[93�2� &O��%��*@G
_Dk�����Ϛ����+�)b��*��QM-~����:F�CF~�c��,,7ދ�dۓ&����E�ԭ�̼�9M�:M'	��}C���=n>���2�ǽS�w�� �.*c�{E͈�10t ����+�'!���Л�
zO���Qx\'��!���l:C�>D��gz������BC�e�_h��Y�n$x��]���"�m��C+��ɪ����4LM�AdV9h����Dr��)��j�U4Ԓ{.>e��V�-��ѣn@`��:#���1+�QJluw��+dp4�vX�{A���B+]t�Zިw������"�����=�ЦL
[�%��:�f��D��pxM��� |��J�(&�_*�j1��zθ^!��NR����Ǜ��>ѯȏ��Ό��������>�x�[G�,�=2����דv�u� �l�p0HJ�|)�%;4���Z\ڟ�e9���xV'JY�����q��ㆱti�b��)�p��O��º��EVɏ������_eÍs\8y���^��6�Y�w�2�0�DU��V�& _xL�k���$u��eAA@p]�.����Ì�O��ґ�橺Y\4+���[�)p����/kU�	|W��w-[a�\TH|O.��hc(�"$	�f(��P+�d�z2)��+jHr6�A\	Gw�S�*1��_��+�&>�BFJ~xEd���y	��j�7ek��Qb�*�����({����l��R���́༣��f���cE�������J_���:xD���	sL��g�``H�W�r`��f�Ö!��Q���}��` �h�,�Z�`ˁ�p�8@T���D��E���O���0��@&��G��͑��Ȩ^Z��B�5l���"ǈW	M	ٵ�
t��A"B�ت���QJ��A�d�����ϸ���H����k�I0���?���(q���.l9�n�7z��;:`���lң�=tH#��͚��ǀ��;����<)vfr~w��%��B)W�	�	[��G��	�j��m2�ۚ�l-��I��_A:p����-�J�����3ڄ�(˗�p9r�>̪�s�KeJ aC��Ŭ������<�a�H;�&�>:�)��+VDT��~0SfRĄ���kS�NK�t1����2��Hv�w^H��/6�:��O���ug8����;^2v����J&B�G�����#Y����\g��0��k�8�|��.3lU�@D�@-�-�!#�e]��m{B몭K ;�Ǥ�����=�3Sk�����N��v_�b	��:Y�RƔDλNSO�F&71NP)ZRϊ�����hpX���,��nr�V��j7�U��P��~܅W�6
 A��#���D�,�~vfdV�rmt.��	�������Cq��qN�Joު�|���R�[��1��(��7r���ټ�*���Jⱔl�ic���B�����||C��S��!~�O�%Gq�<���p�W�?� e����L���U�t���d]2;�a��M�p	@
c�A��@�jVì���m_����u`t����`��ho��985}2V/.8��r�I�<[$⯤h��R�{���̯PЗCq�;�N������.��D�i�c�v�V�YFq��QS\��06Th3���%wt��M��0C��H��t|�Mf~�U~�.;]�9� �[$n�߱�XfR���:1�� �]�h�u���K
�q�w��XS�.���L'�R;^�=��ٻ�a���j��<�p�T#N)'���Ǌ��`pa�Ky�+b��)0s��{�s���(Ǔ�M�׊Y��O<.�t���q�φ�q���52�܆{ո�=ѬT�	��SO���3���S�����&M�E��hr揃)�U$�d�t(�%*t%&���@�y�A�PAPUz3HɡoX�� ��S����, �\�_b����%�	btfi��e�7����ˬ7_B/��M�i;��̭�h�X���g��F�.���*� dPzo�@���U)sC�U�QW����O9������c�@ ���
�������"Z=RuO�����tV���g�����œ�Z�;�`{�SF3��㓓`F|$�G"v��.�
�������6�s�=�{�a���>�MH<�d���%~6�!4@�6h��q]V��tL�I�	�U�?��M���L/�y��/\��!����z [ڥ�x���w	7��Cq�ɱ��"�[Kp���	�y���:h�u&9{�e�ͫ��-J�ڿ{EI��8y�U�u0�6����C�aX���ϕ �-W��DYE��xJ�� t�kSk�W��@�	hH��?CP����6�l�I�	|iPM��A�>���X�}�o�R��LK \`ٝB}6�{#1׻�E��{,�1��#'Rz���b��(��qR��XA��ښ���=Y
��0��-�GYd���m��ТF�-�o���2Ό���w���9K�IC�.HZ^��&�j�p�t���n�P��B�BV{Yf��	+�VO�qw��5�bʅ/'�9��urA˄D��孟�dr�9��"�#]cav���Xs��|?���ty���U6x�O��'Q�crI̧�����G�q芴�^1��4�6޶Y�;��$H�=��$d��v��Z�@�D�&�xg���^#��1�l���Qy���!<ə����T�eA�Q{ �_`�����:ѻ]�^2x�7p�`���������#�5�r^�5]U�_6M�������UB��3�o��w�����zO��d
�p�J��'� я3&�G���j�Y���_��œ�U�!>A���L��FL��B�#���pN,���b���DA��2�����6N��sN؊Aպe�����U�4[@���κ�j��b�/��i�fp9��qdh�N0"6l*x�i��A/q�!1cv|����g�j��*�)�^�x�j��aG�$#R��..g8I��5P_{��Xq���Ɯ]��4 u(·���p���Px���!q�:S<,}��o��C �����U�{A�I]3Y,��}|e�O"���H����R�?�� Ne8�Z�NN��������:gw��~��1�y��p�������[]�g���`�כk�����y�(���"{�<�a0}��e4�&A�����;�Qc>���R$oÔc�f�����@���ۄ~7�&m�=�z^���3���P
A"��?�?�IRW�<`�J0:�bTɻ��[�K�*@�5��]$;�|>Y*oZ�1�[?Cr��AE_�E��s����E��W�ģ��ܾ����}�Ж��H����q�M��]����x�m-�"%���V@X�m�Vo�	c�?5jցU�'=���~a�Sڊ��Gw����M�婔Qt�����8�t�e+���Ҁ�En�.��\9�?�q�J�}�V1(���H���V��5�%��2$A��jD��rz,}ٖ��j�w�v�%��d<%j@�3�~�p�/���V���C���k��=�;�<�w*��)��L�c`�����-��HX��+�)����PB�)�o�M�	(�o��(��:�ԗvA��^��Bv�B�\@�/=xE�><�)Q	X�.s1���%�ehziIa���P���;��2M�QG��5�T���@s��B�@���3���`ΠF΀(i�s�8dN������B6��j���]D?S����Z�a@N%T]��M̓p:S���_	(zSŃ��8�TaG�!�{���W���i#������r�/q��]m��G�����\JصoALg�|U�yu�hc����/_-�~J��kdh��� ?7&Қ�_
�EQ|�������1!�ό+8�v�&�y��=�Ĭ55[��5G�&!<N������|�,Q��