XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���*���vYn��̲C`���]��S%.�Y�D���o�������=����n�f�M�Ԟt���� �e� ?��Ilsʕ���4�b�(�&��"��·@�(��?la�w��o�<I��KבWJ,ܙ�S�=m2�5s�Æ��#�o}_��E%�z��1�u���gWZܚ�$|u���s��л+G ������*�U�V��p�����2o�H8M���c�
�$W9]eQu��t�ᨪ�3��]�!S�U��3-*�F��2�s�"be�\<<�q��p8ɘ��c�]Ǆ._�*����^���<m!�����X��đt�2\�7o��~N����ۤnQ�ak�A��4XS��^P7|49�%��3G
�W��?.��z�Zc3|��Ӵ_�U4G�����j���=G&Hډu
�@��My��_p)<�nRw9�w��s��{���U�-���2o�L��I�'�_�i���ܲ��]'�e���H1���!�_8Ct/E�B��0��,Rf@�`�+uGb�V��L�L7{F��Z��������=w�(=�T3(�nh$�U3 ��=�)f���Y�"!�晨�7����;���9��9���\���!б�*/Bu��I�"�C�3KGKw:�3X(֓#�i轡���<�?4p�Ms�v�e��d�O�ہ�n�W���dAѼ&�u�w��������<f������ջ~�;e�s��N� �4Vt��W��5��e��E�[���C�!)�hXlxVHYEB    1eda     880����q6��Q6��=�vXD�l#!굢|�R�ܸ[����4���2��q˭C.������A0��-RJ��au�$�`6��p�0D*���AɴB>��GZ�+���ܐ�G��絹�T�,��Idɠ�~E�U7�3�#�\�`�>��p����D0uS���)�id]"���&8S���VO��]���C��O
�:�#e������T�$Ƹ�2��b��9��	��`HY,tC7:d��Dŭ�ˈ��5���<��+\E�jfIK�����I
���j�	���^G�/��¾�)�|-ӈ��=v\��{����C�.��&AV3��7�� ��j ��^�����(��~S�1Om��x˹�.U3�$!IcK����$B�7I�?r�zx)6Ъg��3Ҟ ��ѧA�O��:��"4!JK_M3\�GQ;�����"d�����ا�F��%�cL$��j����N�_�꩔�p��W�?�u�#|����mv�/ق?܈��I�zf�S��=[us�"��I�+w�R�\o��v�4n��:��~A#�J��]l*������e�WSKD��0
��ʮo�)�Z�F��R(^x;0 S�o�VHXވ��� \�H8�&a��f��Y�� ��7O.丷fW���B�p��9�Ќ��,�ڜN�W`��ؑ�[��Κ�k���-�/�a�t|�b�←����ڽViְ�͕icD_z�s���`n��{�g=����~��prl؅+�!���w񪖽&l���ƴ�ן��ۄA���)��W��k����!l3���go�@��'#���P�B=k�)���"%��Ԁ?
L����(n��<����a�&Ľþry�O*̓�U6�����4:��W�M���[����� �trikƖ�-�s3�7|���k�㻚h6�kB.EQ]�)"��Sh\��L��A��h�D2��d����9��s7�j1B[���^-�Gr����}q����a���$���_�T�)M4�Γ��S�2X
c����:�����Xb�B��?��`3�n��2��'���]�������25�'�$��=���W�b�=�G)�������B�s0CG;糋v
���:�(�,�o^�|�K�&ޕ��H�tP�r�)=�"gk)�tb����Z�= �dʸ�Ϝ yl��7cN�7��2��y��L��( �6ig��:0��D������LML:�ޡ����
�By���(�ۄ<6�$X���3P���z��>A�;���RI�/�h�v�|��$A���[е^
�C�5�02�`���u�x��������\l��941�}H�m����m\�^R�n��a_�ra��Q�&Qʘ����R�}�TJPڂ�����V���xe������u�J5'/�o\ˏ�'��:OoEo��mbLv�V=ܼ��TOJn�A��D���Q��S:\���l{<,o��������j�)֢�
nD89r�Q��i�W��L%i�8Y�t��������x�t*��]ʔ���Y4z�vH$/�Nu?c��`���𷚉I�����D]��
ͭ���&����S#��QT�ދcl�R6/BoMU�F&�Ln�� �Cj����s��D�	�i��NU ?���P�v��G��=�$jʵ5(ʸ�06�EZ�(sNZ�
"K���,+��p-���љ:�䶰� Ó������v)F�,�R$���'j3��;�M������o�zՖ�f��m�墵th��	Ն2t�������A[*�����:��'ڠ��9�����ʾ��5v:>�!���N����V h<��=
}�����OF��gR��
�����y��"+�R*��|M��жNF�bj�n�t_@!���y�� ��W�ْV���dsL��ru�Ƭ���_��͌��<��u�W��|4g�x6y�Y�%���5���[7&/���OO(t�?��~|�������z�2��ج�s0X�㽞*Ol%��}�[#���
Ó�=��-	�5՘x8���#=O��Gz+�:�C�J6G�����X�����V�A�}�>�1`5�,�%=S+�Ԍ�=��o),!}�.(�����t!����jN�
��H��"H�͡�W�h�k�y� >I�F