XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��AQ�(���a��:��O�����פp �ہF
�;��e#
�QU�1���~c3�ؤYLn����/�~KR2j;K�p�XhU��;7ݍ���\bW�9b�%��[Ӟ�t�9P���`٘Vi>�'���_��c��>���6�B�{O��FZ̴hb>��HXb�#����)pRHНU�3-I�E`����]*�Ⓢj�c�q5�E���� ����r㜁����g�͈��ʶ���B�V%�b��@4�2�S�=���\=��S�[��BjA$�bLj�4"81<��P��xQB����<�U�r��r<z�+�I�H��`.O7*n@ON���!_���ds���5 u���h��}]�� ?�\ u�g��ek��8�К$�Q�j��pp��u�K%Uj�~cs�w��a�h}[r�@g��|��N��-S�t�f��q�z�����9���3b�Kw�i|xߢ�k���"'���I}�}`�l��~�=6[�Lw4TPq�ΛP�������s�Hgh�pHr$E�-rf�=����Yш��
��`&�n�?S�M��k�JK���렼-DUq�$�� ��'A�_fO�f��adKC4�w�G�Wn��l�c�~�!�L��%	B޾�׮�0	�>��V~r8q�>��U��HpM��T�'���|o$�t�����$s�L�	k7���׈����:L9q"�a z\�E
���1Eԧ��2x���<kG:�f\)k����Z�k�K5���p��2�����'\!�A�XlxVHYEB    1a2b     8f0;����Ux��������r����$�0S��������dr�\���A�n���ͯ�Z$�jI� �B����^B`�q��^�U�s<`q�@Y��̠&Nh�i��҅q8����j\>J>堪<	5s��a�N��P��e��ߊM8K��	��-Tb�C�W!�,&�)
	%�;�Ӵ�i�twk���~���h�P֪�
������]�����V���B��u>`�թ��HF'@�N�4�)�{�/�@����V��i�<�ZAY�]3��lֈ�)?��R�*�ۏ�Y/~��!��_��Z3�e�����-�Nm����4p�A�]}�d�q"�PH�f��t��[�e��z����Gێ��KqZ4�As̰P����߅EG���ƸG{7m�h�kI��d>x�
���Z���i�`������gi���⪽�L�'~�n����b]�-�L���Eju���1]����(T�"�!�ơ���<�[؟�c��aF��L4b��B����71Mk�0<� 6>�4�o�|U�㰯Z���  8e$�#��|_n/�o���Q�l�q��}�&��P�<����I�!���(��\�����D�g�f��p+���|���3j7�8@��ERݤ����#�7�ʠ��s/y����q>�V)]@���Ն��C�*Q<���
/;K4�`_pD��Ɔ��-Ќ;0P��9��WJ^bY8'�R?ܒ�E�n��q?BAM%S����˟��5����ǂ8a%/Kă��M�ڈ׹�������o�n&z٨iw�_��ǧ/ވ�c�V\�=<��ژ��^�7'�Հ��C4�Ï{� ��W]�@�V�_����d
�"�Y�)�D>!Ir��� �����pњ~�C���ðm�8�O,}	SW:�ƻ��$���w>�[r� ���͏t�젳Q8�ۼ���y���O��җ�:��{�)<|i�=��~2��hJ\��*^1�Q�*���H��	q1y��{��"�}�U�(�|@�U�	�3��xĴ�	��yͳt��k�����2�����9jjY�Q[����l�Y�Vk6y�-zbOS#���h"�ƙ)p ����̝,�#|#
VCUJ���$���b'y�L�EW7�+�3va��e�\;��Z���
�1�{��VȮ.S�q����d.��a��m�R�RDRB��,^��9�y8v�i����#�ʨ��/W@�w�
L�u���"[� ��'T�"�Q��dq�DX�`�0�ۢz��||�-�D���K56p�E/�rN�@��"	��CH�jڌ��S����#�i�ݣ?[2�UV�_}jύ��D�!��Jg��X+]��{܄��aH�%�s��L;!�וG���HO~��:���-A꥔�����s���� �!�ϭ2=哐����3�����Y�M�D�)�ُ,�Ի���|�y&���:�!J�S���������Q�i�R�!����C|.^D�2*ie������M �D�Ml����ì����S����z��kU>srN-�j����7������~��;��(oǢ=���x7O�B�Y��,��fOHŪ�gk����U��[�"�O&]�'`�D�z׉-�#}d��*$Ӌ-��\��N��ł��\뷘W2Р�a�Vl��lF�kB�/�&sr�BL���Ŗ��R/�VMy~lHX䐾�$�7�ꈥ���m��/{3)���<탍�u�!�2#aiW��~�P�����m��
��˖�٪O_ӳ�����NZÍ���q�IS����ħ=��ɬO��%�	RUꭩԓ;�h�Lb�[�1�����8�=�b�+����_����жeA))��67à�
��uZ�A ����j�j�q�Y�����	>�,<�v樇�b�o��L��(;po�ׅtg��x�����$^X��|��`i�@���wB����t4\%:�i�����??���ps\�F���L��5����
S��4ހ����v;_�K�y��\����*S�j
J�DpM�z�搪��L���+�-�O��a�Y��Zp�ծ��6�N4+���L;�d*(���
�3�՟�F��(�	���|rV����;�P��Z�Fl7�����T_U�b����+���.b8��8��L1�J늩�3�֠y���!�K��e$�W�&� �_��Gq�t��U��~�
`�@���K3 Rė-��q"�WH��J����Y��D�A���H�p�_�[-2�