XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��[90I_�:\��O�$�+wө1)G��N�3�.a-�%��F
&�d�_�o�0��Y���Cd+VpmU�]��K����Zθ�s�=����G)&(��M�Z[k�Y�����ǻ@�wr�)�[��/V�sI���V��Az:(C�΂to$P{[��֮~-A�:2�I̋�����C͓\^�)����?$*>ѻ�/,y�i�,Q�`sς����L=����͗�L��H�k����@��P/ Quzз��#�Dd�x`��?��]"��{U�]qO"j�g.l%����)�$n8{?�q*��b��X�� ��; `�R��t�|K;�⁐m��h��hWS�GP���<,:m���!�/�he�4w χ�W��L�����6��x�
�A�uB��S�����[Z�FV�Q��q���	0<nN7V�:��׺IW��B�&@�?�)�"�� P�`�����_���cDD��I� �o�`�j����6����oDe��]�M�M��_���԰�N�]U�t�h 8�^K�j(����ա%#����7�sTх�X3ݤ��0	�s�Խ1���,�/�.�M�y$��T��bU�l~���R�}�#�ߩZJ7�"T�G��Ӿ~%�3�����%���IڡO^�͏�m<��[碟���-�|�~��r��]z����~�n�����sJ��<`���^��Q��1��v�ݴ�i�n6��3|��R�D�"�4�99�a?��"�^������Jc�3��J�sn:��x�Ec6FXlxVHYEB     f8b     650]�C�<dF~���1kU �L�<d���CD�b1�j
Vަ<ݠÅ�x^Y�J�Fe��+��/ѯ$qn�Y�*:L���u�k']\�eSq�d�Y��,F��YȠ#�)7�9�%�eDh�b{��0�?Y$&�
+s|�Ȣ�Th*�y����.�"]Ҹ��Ԗ�%0�P�5<��3���z�?�'4_8m%�������MuS�_���I-���-�<�0��N�iq� Zí9����]x�N��uhRԾ�����Q�5�&�g��NX��T��C�
�^v`[ߠ�_��վ�]�8�٩�H�}2�J=�"��4^���$1D�5�W������s�����
�#΢�6B��x���n�*�F4�覯��V���h��G�/뫔9/"\��&&킐�)�ݹV��eQ����+?����_��^�ɠ��o�}�����)�A��g��_j8�Vc>8���%@jj(ϛ^ � sc�W��7��A@���u���U���k������	�Sf\�+��~�6@pDs,Ң��,�U���l{�Ol��_�~i�1��o�j؀����B�-���5��ʡavi� �+�Ζ�b+���8�?�y����P�񟁅�g�s�cQ��܃R�}ok8��9���uAn�Ua)1U��T���i�:}��6��R\,���V���dK�)S�c��:���ʻ���˺Wq_Bn�s"�������/���]�(fcH���㬆�+����P�0�EXLY�3��-���b��5�º�",7�A�C3.�F�d���Z�b�}�AL5���ր�w)�����t1g�~�&�dC���brt#p��<v��$�>�~�=+|��p1�ы���z�*�7�����	�h���>�̿���d�纇\����8�.�VA+)�U�����kjʕC�O$�2��k9gV�O�����g�LE���s��{�$s��x[cj��+]*�C���XJ�IjOO5;@h�t�cVG�q0�Q�DW����`I��`6}	Z��kp7���=@�DM�j�(�_��X-�����i!��.��&��	���E��&Ϻ~�<D�8l�z��'|m�?>�$��sc��e�z{�y�Y��jT5Y%�?���SM1��K_�/dWe���˳9 �(��������vc�N�c��FF��\�Ǵ���m����Ƭʘ�/@d�$cgB�� ��WGrr�[�-�t4���
I�8z�4��@\>*�E)�W�)� � f���J��m%�?W�����hzc��ᖮu�/�>�{�EG�t���� �"�Ȱm9�Pt"�<�Ƨj�����n������[�@5f��[��m����t��P&IJ�����L�@��S6�"��W��U\������aޅ��W���-�T�"&� ��q�\��*1�?��%W-�s ����9���Т�a��L��e����(t����e+��%}>=<����/>�o�<�?7�ڬo��s;if�z� ��\:H�s��
o�A	K@S4+ԒvA �~���+NWI5�*U��ςm�k��aj�*^��w�#��׆���*Ϧ��Ս�_@�^E�T)� ����W�.Q3�6G�]��lwu�au9c�h}