XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���t>���܃�R0��&XZ��g��z��u����pU�x/Y�cl� >2 `e�Y�ڠu�\V
b�5��)�;�p��4y��G*�g���u_3
�>���h&AƦ��bp�N%���x�쉜2p�*�seOl1w���qӚF�O�YY�dwX_x,��agh�f�Y�6��E��Ե?�t��i���ɹ���UMsf�,X���,n��Ҧ�����K�Q�I�*�������}���Q\�d�_FOi�ܺ�8z���}��G���n50ޱ�D��)�O����Mg)�~�E��d�cM�EΣ�@�R���I�^&�)dϯƍ��Wl�@�.^o߶i�N�@O��\K�kHΧK.4
J����3�}J���\���?��¬�����28'�z�"*�*��b9�U>���M�����N)��7�
CPZ��Sҧ��n�Vx��a�x�yIK�no����a�ps�p�Nn:K ~�.�<���+���F������u��(�ō݅�_���q#��Q8�W��W���d7�K�b��B���ޙ���(=:���9�/h��	qP*���0]��:a�
9���ɶ�]���Ŏ?;��L�Α��@e5t�R�߆�DN\+C��gS4DX�1T�,�T����pZ������^� �b0��d-0ܾ���V6���@N���-�Wm��0����Ť�?����u��_�J<,kG��p����0�5�������%�0��Q�_ˬ��0p{W��<XlxVHYEB    4c95    1190[�Y�G͑������[6t�QHO����  >��\��o-"Ef{s�A}�uL�\�����SK.���kW�k�0;�����8���c־�>Cro٣e�e��ęu��@k,L5��[�Ǧ��Y'���Ӄɮ�H�LP�y�ϵ����r��
�m^Dg6���5���$D3_$�mŃ*IN�п�WZ�˷}��G���`�j�1��Q��(˅&����s��s�1�o8 ��<�9�vU�8�ܢ*y4E��9NTq���a�+b�M*�;:���to!3� �[9�0�G��M��@�{?9�`�s�����0E������1���=��Ǖ5��2+�pL*
ʤ�V�Y�$.T�	�V#C�zY�d:�5�������I��`F�Ëz�>�c]#�κB\^�=�us!5I�5�)�R�a�G楹ǚ��ĐG��u�tM(rr�g����U��`����NޤJnug�Ae* ��y�`ɞ�W��{x?�>'����*��H��n"��T��0�E�X0��*�j�
��]�7�}���ݵXܩ�S�U�d�3)�`�VT�3��E�Mhb=6�E���9~��'�� ��f)�+;�H��Js���=������z R�A�҉͹}d�kR:�?Oj�K�X8��Kق�HA����ֱQ��l�avlz����ʧ�i�e	UӆT��h��Z)pU�[+/]��OH]�R+���0t��ث^7��0L%���3or+N$���Д��7?s����I�ϧ�_�M3[�O*뒉�ڴD�NM=��_�N���x	J|�_x@��c���
@!���R�)��b �o/�ف%v�%dt�`����	,�x�HF�/��u���)���ϕ���Nhʘ�k�SUg��،yD�0/�rD��1���e�P�@�(�e��8�I�_�ᩢZ�UD�"�l�f�D����n��_��ḳ*���J��x�\��h����v�^���y�h�SYϴ����A?� e���L�k*#��/����8O���3ŷq��\U:���3���"�P�r�� h���� ������+�OD=0��.��q���Y�m*@��)D�VhR��B.0�O�A.	�]}�5	�n!�x��	N�^��D���1z3j}�+�=e�#���]�!�NZ�!��aʷ!�`3�ۂ8����c�Ggd)�D˺��KΘ�lˍ��;2�>���+�����Ȣm`��/��*���g��I_��kf�fn��g9�?��o,?���%`3��Q���
?@P��i�)��%��F��qf������`��@jִ��H�4́̒Y����� [�V�B4��C�*��8ȁ�l�ny�Y�H-?kL	}&ܺ��+g�W݂0|Q/�%�!J@�o�)�f	���ć����d���WSO�v��ݐ�i��s�U�u٠/<����o%��?�(�q��^C ="�4v�$�A��G�Af��&ڛ��I�g�B�܁� ���0�Wu�SՋY�jc�Ҥ�Z���d�D��k}�r�2�I��?���-
�2l����58�J�W�If�EC'l�o�C(��w6<O,��:��V���a�r��Ug�|����κ�v�/^�N�qz�P�s��+�Q�Җ�a�+���($ʝ>����L*;n�����<U��(�E,���#��ND" Y��\�ڑ�P��6\�������Ȋz��p&��à�����`�i��]
�Y/}=Ᏼ�0|?\,O���@����wvIW��{�c����@�d3���-�lޖ��#^�
w����a#�np�j�{�9� �/��D#H���<��,i�Z���I��`$��&�H��2����S���6�!6'�����5EM�i>�h!x;�6fQ�|:�qY��T�7�]��7��O `V5DS�=��\Ք�O�ar|�B��E��{��(IgR�"�'e�ּ��=��K�GF��mR�ŴeyY�}b����p�=��+��~J��{��F ���1@�W	���	a/�t���r�����]���ֶ�n���!��B�E��8UWY��1���@�ʷy�8�+�\���1���T�qz��h'� �f=\�5��������X�>�_z�������=���ؐ�2����񩡑�5e�r9 ���	-�i+%�=�#�a�՛��Z�X���P6-yV8�!p.2MV���.\N�kE�|
?�Z��q�AmR�# �5�����q�s�1���'=Q"���^�(L�[�#z�Ů�E�`F�PW7�EW5�����xE���P�)�5��ػ�ѩz��]654�|A����f0��!'�$^�ra�x�s�����9��ѓ�E�DJ��E�!7 ���75�@=�Z<��厅���8Q̖��mfȢ�g�2١b��v��,�B@f��#N�e�����k�y�p`%�Ҕ`σ�s3ji7�	��<�DPd�}r;$D�=�_`��|���(�����'0v3�OO<0-���������2Ju8~�.c���H�{�.��_͒������%�I�R J�)gp�U��KڙB!�p9>�EXSf3v�'zc�˽S.�B#M��l���l��_�Ԛ��܃�&R�ɢ�̟��������<��0���L�!S�q��x���ς��u��1����ק6v /��{̝�ZI���6|S ���A{��g�,�x�e�w�@F��n�f��y&c���:�@G��*m��<�ޕ���)��&��_�`ɸ��T6�.� �����p��e��H��|��gT��ⳣ$�^h�#���_��~���%N��d�O����f7���eւ^)�81)2(��u��#��1��5[�l��)�Et��!y�Y���8����)��Vo�W�
j����i|��1y����|�Z�m�=h{ �~#�qn�e��c�3GL�3L(I�ƚ�#�2�_\�_����>��뜱���:L&���d���tW�3\%�°c��O�Ff�I�'O�Ta���E����A6j#aj��i.�����w"��e���)`>��w6���i#2%<��j�i��C�i�F�^g?�7�૦b���Ra�[��A�������шc�u��l�{�Zv!��	��e۬�����D���[��J�a�x֞ݵJ�:�����S�y`����š�8T�r�ګ��h����Y=(�\0�$X<!s�t���O��k(Z9��|E]�����J�������ыi�-�����UEA��u<�k�f�����ڇ,��.�pܮ\z�*f8�=I��+�0ގ��r�o�nb��k4�TjoFҟv�)}��?wZ[Ҏ=}�&k�S_�<9uai�pFK�;k�SSn��5fM]:��)������r�`i:�;�qǡ��ѱo�,���Ce��r��U�8H.pJ=4"�o�p(��<��_�%}��s(��c 9W��NJ����3p��.s��ܼ�u���w��#�f���*�+s7Ke���'�X)/� D
���9���Bŏd�	��+J����@w\1o��@�hk��SY���/}.y��$LR�8tL�j���8nH� 6���u�D7����57��asfV��t���̮������s��(�}ʄ���0��G�d�y)ߘ��Z�I�(�F�3�"���f����3at���8<Dk]b`���M4ukXX�є"�c/��a{��c'C��[��b��ꍞ�wvm���l4}V�x]%���N1e�W�~<�ǝ�F^#��I,:V�q�D���9�,���)}oF\"�x�[j�$J#~]����Y��[]ע����k���k�*9>��Jk����B�BYp�"��>|Zv��ϲƨ�H���{X�1�N-��\pz֋/�z_��;|��Rټ=i�=ę�(�T�8��������Z@D��9P�l������*�ٶ���ǽA0`|�#&�{�ڝ��)s�W���r�3��`���*�����O;���9��
N+:�����D�E����i_��/�6چn��@�j���n��Ų�ё�D&c��'����Z�N޾^Q%H����I(�D�D����=��_.j��	����t��b\$z��s����{b*��\"ܲPS�"<�0�:�X�#��)���~ǐ�ڶ0	J�PW�S9��I��\b�W�+h�A��Cs�Բ�R\�ڠ���x���afb�ΗɂCE �p����UUBۦ|�#Q�0�2!�8׉�sN���p���t9�"�ڡY�&ͬVD��'!�Z�El�w�/�rJQ��:��v�G�@�;�;�3n3���b{s�M�<뢥�g^6�!1�� w'�<ɷ�I���+t|��