XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����K�6�ż2�y{;E�yn<�\�Nb+LSn��R�X�s�Y X�5�����1�I��ۖJJ�!��~�f߂���'Tqp�&C�5E�p��1�-�.�߯<�ڎt�F4��`�Ӟ�GH��0�q
P�~��ߙ�g��٤�����,@��G�&/�<|�N���~��v&9�%v�O��|R�o��||���ȸ��� �a�PN���%�=p*��(�>ћ��ě.#-�fm��Ī;n7H����y���A�Xͺ>�Fݞ���#E����s�P����Tm��*ɜ��WѤ�4ll~"�J�$XêN*^t%��Pdr+�@�]gT�c�Nu8S�8��ΰ�nD�.}6�38��d|��v�&�v�a��XT0v.^"�B�rԑ�)Qj����$Yg3�-:T�H��"P��"	�
.\��ӑ�ټ��(Z�����:l1F>W�e��XZe�{5�;Xv�J\��)&��!��|OcMGz�踢ay����(L�k��)0r
��.M8~S,j��x�pM9�F��6�ܝ����x\�����~�%i��zƠ��YQ�Fܗ�7v���Kg
��b*n�%�?�3��Bxſ��t޷�$�b�V����"Px���n���/=�!��D��27?&�P�J���<�}��6���}� ���d���U|M�i�%|{�*@=s���H�
Wb������W���O��T
�9�L���M��aiO�Z��l��q ߊZR��G�1�M9Iע���m���r�O͆�B�l�$TBZPXlxVHYEB    18fe     880ŭ�q2�p�:m�ŸŽ�\�04��J�^�߽ѻ�I�B��>��,rW�C��-ӿ�� n�����:���Ꞗ��Ӷ�u�8��X�Jz@��.i|;��{S�m���iO0�"@���sLnM�a�A%�V�q���cƧZI�O�����@�V���uO��f�yLX�] �W���^�a{�	��$gBq�}�&�|���Y!��.h���o+$�:9�)���VT@�j�5̦�,!�:کA��(�_ӧwv#�5:k���/�3 ײ��ѧ _�_8N�PBÃ鮒K��/|��Ӯ$�%+�^]��w�j�鿸㐛�K7�_8�3|��L��k)�
Tsh��i ��P%�-�W�Qp�zִ%�!�lc1$x_��&���[�����a�A��>��
��c��#B�������G��q�]'H	�lU�1����Y�vR�FV'�YLj_�%�P��IpdE9�m`_w����}�(�Z���oʬ�� ��0;y��XZނ�=i�K�l����$��|o}���3^��# ���I�g}Ϊ1\lH�ü��$��ޥ;?#t�Q
.WZP�o���@����zɬj�ASoH��3��u���?	߈g�m:�.dD�'���ؤ,���b�5<���>Ǎ�M����{>��'�	04n��;��QvZ�B��O��]8�Ʀ���p�r���=A_N0͵�]N����Ճ�M���tvf�����V�j��j.�C i�R��.p�6"V��G�b��ڒydNr ��dAf-��4ʦ��'�q�	�h�m�-�H�8�PqE�*��|��ϕ�O��jy�+�\��[d@2v�H��U���΁?�'�[��$l��(�*��ث9A�'[�^9�21T%�	��77�����#w�(��b�������uZ����=[z=��m�*]�ӏe�H��W�`cA>D�T�9�u\�Ć} �����z�����FI�������tӳ�y6(�Tz����p���Jϒ@����T���8�G��O����sl���e�3jR#y��<�b9�چ~a��Ju4֊x�����������-��s�����{`|�sک}vOK�)1�9N�l���=c�m�H챜͑��4|}��}3Aw\3ŏ�� '�s��<��h��&�woT���ju�'~ƐQ4��GUO�pJ��b"j輟4�}a�dv����nP*g����w=v|�N�v��O�'��z�bt����GY" ��`�y�GJ�@qWV�-��?T��`)�,��JH48��<�3��;4��{�ދ�¥�`�� pm��6��%�I$�u�~��,兺�OH9�t�$�q�Έ�Ρ���;�ā�Dl��v� eǊ#'�N�z��D��g.v�o��j�aO4��_�
S�ƪ���7 �)b�%�r�KWU�9yKg��.��͂�naAGj������x�m�JJ�0��8g��H�b�x�6i���'��Q#�m$��,H��Dq���:_S1~��O�Г��r�)J��E��s&A�{�4�lyd����)�+3��<#��FZF�B��'��Έ҉��Ӝ2LW@��f�U��x#�Y/d�U2�9O�x.s�b��O������	�� ���",?9� ��g_SUױx؋�"p1z����p�	7|l�N�5��t�NKx����(j�÷�+#7=Ð˲	օ��x�*gw����!�.(B��������zAd��K"�WjH�K�Od�!�'�P˫7縔+D)��8�V����D�	��x��|k7�,H�bi���\���Њ�]4�R��~"%��� �t�2v^����N�Vm%�FG��Q��#�6�&F5!�,�w-Ϊ5r@u?�A�ǽ�'�I'�ZFq����wFN��)�N��t	��].^��OZ��1��'Z�Ԅ�.����V�Yz`��Vz����"��;d�?�GR���x� ���t��d����f!C��&@��=�!���pkZ����E���k���1GIW1)@:B����
��.A�#�d�A�Ƽ8�����V����?�@tʹx`��;��m�Gj��+��n�,�sv;�9�����SS\�������4OVX�+-~�WeEkʐo�R1�29C��
�� ����o|���P�1