XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��
�!�N2~�Ӫ5Wy��
 �!��@8�gV�u��"�`�#΅y��2�/��4�D�;��[vw��%xmm4�~=-ga��lQg��O�|9�k|�:ݣ���e3CY���P,��k��2���UCd5�W/^�"u�^������-d$u_Y�,�C���Sv0Q��H:T��ߖ��Z� ����Wv-�W���&AbȞ�#��Ak�,AR��1x�م�Lذr����40��x��)v5JK���mJ�n��TP��7��9_w�͗gB��e,@�b�j��.楛WVsX�3 �x�YC��YC FP��:�hKI�5埈�/�g�����`RPVL�M�d�h�1O!�\�
�F�S���H����?<+j���m��j=��π��2�7o�.2rʵ�p�=3i�/-��h��l�5۸�qIbl�d\kr$�<n���$\A0x[BFN���a�w7}N��Dk�o<w�&����A�aD�������\h"���z��<�Z�i���p�O"V̶}��ݱ��<�L���uif��᪽�8�C����Rb0 bI���8{6��$A��9t?{ ��?��!J{V?!JZX���w�(Q��4h�P���ƪ��2ǅ<��0@��L��E�mPbK�Uv�f����7�h��㖭��_0�8�;�j�w�Ŭ9�1�ؕ���V���?`��l��|'�[�`���^m�9fL����Rg����ՆZ����S��L�5ׯ�#��l��Cr��A��`�>��[@
�r7FXlxVHYEB    1231     7c0��=HWu;��ݰ*�P�вF$���|�V���$ҵkO����#���;�e�n*�8�5a�7R!��ɤ�O��Xc��2�m�q�/F�S|�&(P�\I���='����6��Y��v���1�	X�љ�/d��"9t&����L�h�B3%�*�,��H��tZ+�u������B>�{�rQ'e�a�a%���aCH��[�
f0B��+ x����9�Ą
����?��N�V/UF�ґ��P���Jn��2�t�L��� ,�@lŗ%f�;v݇Mq�)L5��asֺ{q���E�y�y��-�]tՑ���$gQd��Z��m�Vm����U�A?9A�O2���]���Q�6;�����}!�DnQ���iei�h��l�C(��G��.#�l�LL����@�]8�ޮkr�u.�M0o�Ol�}ui�����P��:yL��t�Ijs7W��a�kjH!t�.
Q�ODf1�t�R���Z"	GiU��(�	�u��LӇ��)�у�%<�Z��{�Ȳ���?>�c�ȬW��z�L
��?hȳ������K��O��AwAn���(��lJh�j` ��w�5M��{��(M^u�X�H�l|�c@����K(�O0��#�y]k��a���" U�p�p��FN7���&K�Y9�H���=��=��7L�:|��5��r��$@})A�<�Ul$�5ׇp-*�k�7l�Ym(�ü]U*-^k\W={z�+�:� �l������f������V+��Z��q�2'�ޒZ�|JO��Q�q��DO�~L���!�s���|l��H��[�u��X|���5�v�^���㪛�-m4��W]I�<Vn`���H����Yf9_�2=����Q���D�j�����)g��`�����ZO}�|�r�w�`�������l��4�~�D���g'�;�=�q��9��Tl���#��f���]��%��."T��c|�%r�l�j?B��$��lc)"�Ķ�����I��(4������	�����װEHQc&h����w2J�\fV�߼�#���[Xn��ư�I:�) d����.* �GK�D��϶��ޜU �]��p[�*4v��;�'̍��Qf��X�L���d�'I��������D��w$�_y:���? �s�؁�Y))j?�v-;Ŕ�/�ފ0��9�v�Ha
�x�i"d8L�QP��|7F�jA�k����O1�{�b������M��`�g�"v�4���������!D%��GYHe� or��2�z��E�99]ɺ3�,��^ KA���,҂��~���o�U��7�O�(���MNT_5���Pf��Kk�C7��;�L�}x2��x=�P�����0�f2�M�^D��n}� s���C}V�E5�&������D�x =V���O���e�..�}�N��7�{�G T.�(V�����Q˰�����j�r��0�kDN�ƀ�Cj-�e�Z��a(�a�/��z��?��)5�K�r'Qf�y���0���Q�WrU��Sb���� h��Z����@��<�)ĭ��><�ϖZ����JO�=�ƹ7a�)�Al�>�7�F?*�?��#\���+Dwû��C��v�F�qF��n,�4��ͦ� &w�!>�񷆲���𞸾�nD{�};d����#�7r5�݇mM��	��i�r(���Q� �gٸ�Vt�i��Uk�{׊^1�"����j��)����>��A�Gmf���.7���o�;���t�ˁ�D�8��_����B���Rؓ	D�Q�'6^���#��c�N�����H�JT��ԗ5����,G#S�ҍ&��KkYs�ڶp�v�GgbZi��I:f?��~}���l�b˴D�U���q�("� �t������.��7U