XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��eqAI��z�_�_���#�Ki��c�d�$/Q��LI?{����Z*���)�,��}��F��Z��I���r��3%�"�b������I/��݊����Gy���^���p؇�;��J�+�O^8�Epaݵ��L^�.�y���2��oZ�x��kT�{���zdA�g.B>}~#w��[��H콣}��X��,𴉅���o)u��E�>2K�~�Y*v +��Y3��w���	a@�yܽ� �+��.��%�\t��5s!�\?E��W�(i�:1t�8.���/A���c���jV��΋�����c ����f���=+C���N��M���+������m|5CD�r�V�·��7��0�)�[�V�Fޫ�"&&�#�=�Y��엶y���Zu?A��_�:��Ǖ"mtGy��=��<Я�TY�Q&ؚɋ��%��)mќ�Q����=��h�HYo����+�|U��5@x��� ����EO����D ��*A�TSb���ޥK�5���J"dM��ϴ0��O�F�Hʼ���*T�
���ǈO�r9xxMMj��}<�|T����
!�F������%vK�q��\�+Ã��v
�1��z�(5���@��M�eι+�}�~��댖 F�+���n�s�i�M�dQR�?|�Kگ烴��R�`>Hou�6}��u���a��G@����p5*j��\-:Ly d��¹�)N���sE5\�Ѷ(�Sp=�W�|�ԫ��U3Gˤ�Zn�UVIKL��U-��P�_�XlxVHYEB    7a7e    1af0P���mVn�l?!��Ԓ9�����>d����Pz��x]�qY��y���K�Q�uy�*��T��bЮ��q,�����]IV��N
'&�A�,DG66^jY�F��uhh�:����f�8��:���;����kb�)G2�5����?��^`����H�����/��[���]�ή�����a8�/�Ո�caS�=�k����,Oh���q[�C�z��eF�l�fX$$5��+)��x�l�F��Z#x%6�F�wKx�>5}Jl*n��\�e��E���DDƋ���W�7�|���s�d����EcC5�Y\��s�,ȅ<��p9p�r���]h��AVà��+|93
�xe����L��J�G8��ô'�nJ �́�
����xnj�`H��ՠ�,����l1Ů�9h��xJ�S�-�Qc�*I�r���/+���;^��d�S
 �P=P�����l�ɽ~��D���H���G�3u���l�}F|ir�m�9�w����!�<X:�ɩ����#^�fi�>`ѯԗ��>���?%�̜h)&�ށ���Lw�-���]k%�-FM����s�B2��D3������o���u�^݅��fLnT�ꗣl'z�,:��x����t�&#��?���y>�}��HG�I��`9�L�>C����VM��x��3��2��ک�$�K�Oq3�*��R�<��r�Dmʯ�8"��0e�Ta����DA�s��@��·�9��%��=�\�I_�B�[�t`��'r��S���[�i|��K@y?~�o�7XVepY��2�"_'�7�."br�:�JB�07e�$�j����]D�OѺn��J�N�ky���Bߌn=�{i��G����}�S��N�6�N�&p ���`%��1퀟-�"A�=J��>��i�>����\��	�,�a"T
'�����UK�q��U���Y8���m��ʢtζ���Ź�=jI�������e=F���)�c#�=:�y:k��{��J� �0�S,X�)V�5%�'@�R���s�~����=�i1'i�3w¾�⊾g��!�j�$�Xm�rU��h�ms�˥��v���5�)A~�������7�kv�޵
(�j��͊f�#��bũ��1g�'0p>�*e,�o�N��9���A�p�*	,H��j�lC{��E� �]_,h9f�̍xªkK�Z���u�ER���UxSn*��	��x�]8]\�{?��y�NMd>Wּ-(��'銛��	���{�s9��b�������;5>��4O�u%�L��3�{뇓AHo96�&x�'�	�~3N�����T���,X�؄�W�~�s���q�&� 8�Ű|����g>Uu�o�D���>j�%H[��5���XdE���k���PvƿRK~�𢖦s��0ui#�c���&XXVQ4�`���	�K�o8�md�7D��� ��>�2�'�b��D��I7L���Y�o�I~[�=��\�;�`4)�B��A���rTM���"I���}��a��Z$�@�e#
�.c��,a��?�$+�[4=ŠÄy٦|���y!����q�=����tاA��������*9������rf�AS��}{s�+���p:�ݵ�������0�J0��b�����Kq0�x���B	������O#�u$"����Գb�zyx���*�ۛ����Ynȟ舯;Ƃ���0N`���u�{��xސ���Dݫ�~����P���'jJ��u�.p��/�Ϝ�湿�6��#G�<J�b�E�'�{�j�d�'+���k�16���Q�$��_�ފ�;):Q!f~Xގ�b����i*2��^0�~��	��I��Y��{s�
�(C�O�}��Z���|�<�R���3*\�	���jWl�gsmｳ����UC AR���Op��h��J	��,�S���!��;Pnw���ɷ>Ֆ��T�� ��,T�Q5q0�fns�kSh��|��='�V��r�ݭ���>�{����U7����c�2}s��,F�VƷ3`�ز�m��}(e},���:R������bC㺍��n�Ѧ��VKd�&&<Wkn���+D��v/�%2�dУ!��A�z"������.����~�Dr��agxj⻿jYB�Z@�n�W���������<�^�|�GuN��,W���L��ۧ���(��%a��-�vZh���^9���B�0��f�����Mc+�v!O� �-b�
���ڠ@�AP��i�w
=�Ei�\�ps�1M�`�/mײ��A�Fu��č]��bw[��-���K�{��y5��g+��Z�l3�寲r����v]��t~�>�	f�8E�)
�L-��`I ��%�����e��� �U��9����[�瓬,5��
�� =��'�=q�#��R�*�`K�~�
��4g*�B]�H�D;w�|�����e�a��#��o���{��)����-7���L}(���|����;Y�1�c5G�-6������� ��ɞ�Yf1�tS� �h����!���d�{�������w(�]ô�k�*�z>��Z��[�,�7���px!�<��I�bh� _m&�������M����yF���kCsKV���T�I��t������.�J�L�O�O�f.@�L��7�p<캱8�6�Q����=Nh��!VG)M�*�N�)@��6fS�b�ǚ$���x��_m�L���ۑ�����[�P�o2Τ����Lqb��	���@�,>�*�E�V�TIމ&��$0A̯Y,��zM%����i��]z��5�oH�=��|A�T��dHa/���~}�T����kb����Rb��A���O ���,g�>�Y)��hf(��N�Ww��:(Fn�W��d0f\�`[B������`(�[�B�}�$�D�J|ƅ�qƯ?+m���T�[�.���B'���A3!��o	�>=���X3���(�!p~ph]S\��n.K�u�U�C[R���MHh� t,n�_�m�0����:�Q2�n�J?.nD��IOޯ��E��B�p�䎹4qN-0L�c�p�O_����6b�Na��'ZdF�7����x�m�
g����� ���_6�σ�h�ɮ�+���m��:���d����[Z�M�Q�s�fIc�����Ǜ�U:�B����N���f*��i�p/g��Z�8��������x�B�ī��7b�kj�b�����p~�o���T�+aT��j[�$�V�����g��Cw�3 9�&3*x#��3g�:�V�����&�����2�Q�=o�g_:�R�[V�t�ZmfJ�*H3�4����v0~w�m�f���bG4�?]��[�F����R����Y��A)&y��cа��\ؚ\����s�y����a~f1뜋��&U���%{�:3C��Ģ�"_P�%�3�ǈ~6�� |��_��:e�[�2`���e���=�Nꝰ;Vjŝ�\!H3��ܬ��XMY�'  ���{�7:J���_���c�S=dAt���_�e�|���-�4��c6���ܾ���nMXi�O>ꗰ�R+��kYOi-�G�ǢR"��q2�/"��T�_�@��Uz�GA�~̕�0�1�;`r����#�zi������k�I��Ww{ �3u
X��&���ĺ�������濿�)̣�Gؐ���d4j�/���v�e���T�����uq��z���N�&��xϜ��2D���������+v��%���F�V�4F��3j,xs:o��.ӝ��[E.Eة3��;9Ɋ�ł�6���
_gs?���?s�>�SG {]ȟۢTop3�O[^�7ae��@�>Cp�Ԝ�ߙ���=+V��M�X�\�o�#�y�A<�c�2�@M���ei��s��Ā�s���ʡ8�R��Km�SS�>�	�ʶ�RF+� ��.�~)Z5���Z�oY�V�O�I#^@o�f>��q�C�.)��D#90P���j��=��:�L��B�o����H�DS$rE�	d�>9�4�������Hb^P���E�w�J���C2G����.ve�$�R�����ؗ����u�%��_��V�'<�/��Fie
�x�&}qx��� ���t�w���Ch:�����=�F��W��-en3���D;KG��oΊm��Ο����z�io��$��E�!�ׄ��5?/��e���R�����@*�ў����}]9)�W�c-"	"���8B?��{+�Np��GF��*i%!��hS͔P���J�&��M��
8��݋Hpj�g�42r�����In:��P��1�������=���M#��k�&�wOY��HZ陡��ȶ��z��ɬ��� t��pr�)�p�N鱎��@X��-����U{���r����sS�{5}�g���gѲ��c��1�Uzd	��9�qg�: /?7T��NA�	��os?ۏ%`�ɌC2cm�A����<ǌ:h�!dv�.,��
�q���πI0-}�U�il
NIA����W��J�yC��@<"�@+Q���x�Q	��Ww�\��vOli="���fi��T�7�'�`���f�G�FK�9��������4�ڱ0/ըrŖT:7���,���}i�LÞAb��=�Z�2|s�����|�T���l��_v{tHM�#�8SF��N�Yͫ���]DK�H�c�=^
�6��x�X�O��� `����Yxxɤ���L����,����a-�?�$���̲�︙�{���q�T)��N��Yp�
[�Hթ@�	*u�ݸ���d��(Ƈ2�uHe��BV�� I���C7>����i�Mh�a�r������?���d�`�b��̎�=\#�8�K�UL���c#x?6ں�����M:
K��I���w�K����/yIxN�78�V3�P�p�긺g�yZV�md���fq�S>�Ã(Hx����rT�����)(f�P��e
q��	on�|�P5C�'O��B�uҊj�.�ɼ�=�x�]�!L���>S��	] Q���x����>��3��9�)jU�1���nZT����7���� \��&��pUH'I@��84*a^�t���C���A4r�����:����9�@��}��K�9is��n�8m�׹�(�%��*
I�H�6Y�
H8�_ܖ~7���G�Si@�@��̣aS<
(���\˔��7IU?��5H���ܞ6Eۨ+~��/B�V�����#�:t�lNs0�4���V��e���̹z1����Z�߽���I͖	Pn��sP�fU��>�y���l�ԛ���=ǃO���,n���h�J����67�$�����o_����  ��B�ުv��:3S[`>���{���ź������_��](8���V@O���������1o�J9���tQjY�1տ�Ye��3>^@�,�I� ^H��w�%{�-λ8��Z�T���'O�Z\�ɑ_�XxNR]�T��K�}6�D�����Q�^�*�Hqv���$�0U���s]�:@Fg��SM���r��ڬy�x��g�]1��b;���@թO�RIM��A>�4��+�9������a{C��6Da1WZ���\�,`!�����0� �F��	S����䰞��Lk��ƇIϛC����-�������)jԴ�jT4���J��W$�j�H^F��	��]�E�^l��m!��;a��S�n�1V�U�P�7�&c�C�Δ;U�G�l0�X��AԊ��:nŶǲ��RI���-�����a�y6�TͣK�Á*�a{��Ti�
(��z�]Op��J��bq����r�)�����t>��:��9�>(�	a�^��G�f�x����l��.�[=��@d�:]��`�>�M��AҪ&��-B�'����Ofc+��Kp��x�j��R�Og��V��
�`]EW ��Ǉ�B X,��� {B�j�ĎE/@1��!�\`R6��2 ���!%�s�nK:+��2]���Ƣ�n�(��>��L@H��s��h����O�z;��w1��2�:�ߕ���UU�&5646=w�O�OX�!�ໍ��"�AEf����#h2�3�ا����� �{�G��Q��e�䶭�;&}�z�O��0N"f�濛V��H�~���i��p��J��dzhn4ڰ׷�=�TKǊ]���s�C��������[�1dLޡ�H��"���}�)r�ؿ89��T2<���e��k�[v��`�|����fx_T.�SŅ}�Ԧ��hw��H�Թ帝J�E���T�sd*ђ7U��D�r}��{�ƭ���J�A��r�Ю.f��T���4��M�ʨ�^�M�w�����2�!x���U�8`�,hi24��ˇ��/D9L�#��K��"�����.0���>Y�x_�����;΁Uk	>l�_h�4�P�!�(���K1�_�ѾћhΕ4�`08���r��z���{�@�r������ʟ��c���@�G��䦼�n�{$���6u,��F^���P��K� �4����:wB�����2���,�8�L�1ɛE?Jq�+���S>�Z��O$�Y�Q��Ǥ#��,Ǥ�T@C+u�/��޿}�,4�U���άQ+I����8�P-�P������Wj�j���sfRK�NT`j���*Z}�;�������������c�U�����N�J���R;�.0������r��gr ��G���Om��B��c(�kc�m��:$