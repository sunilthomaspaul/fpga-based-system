XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��g^�QP��Lm�#���0�d��AV��9�ܖ��'�y���@u�;��.���;�EF�މ�t���EQ���1)���ѹ��md�=Us7�N�|�j��nF�94UT��sH��NĖh�/�e�㄄3��;�[�\���~\�~�/��߮B�V<��s�wbq���N��\T�T9A�M�|t�ͥ�;C�Z��wl����-Y���L"D\]Ѻ G���`pݓ��4��z���G���;�_L����M��>��0?Ƣ�I�{4П�le�b�K�4���,��#@z���֚�}�6+S!&� c�O\	V�j�`�9߅
��e���pE��;��5#�������7���. "��r?�jF0�6�.�D^��_�L����U5����K$��A/-~��� 2Z��ǺUl�����T�����CǅZ{g����ȯV3�:�ҷ�'_�o?���;�o𤿴!0�S��E)�^���VZ�6�=�>,��3Z4
�g�"�R�sG.'�O�N;�O�����{�ιG��;��$�'�����̅(ƛ��+PsEy�t1*��?�ܵ�� 0���7�3<-=�׭�@w�]%3yw؈��a�z���Ȃ.��Osd�K'�i�:n�����x�ZL�O�b�Y|t�����
�s�X��S%JѢ6jb���H�7��'4���h)����������4V���s��Ybc��D�h�� z��m���!9�d+��'��d���b,��@��s����XlxVHYEB    18fe     880+��Y���� ���z��|Y+V�׾��q^u9"%��w��u�huX*q�jڇe���sFlM�qR�6��T��&�Y��#�X���{gMKW.�D2��ݜ�xz]���S��z>�BG��I=a�$.�I^j���w�M:�&�.��\���T2幯�O��cf�q)���u�C;'��? ��<	a�ZA^��\5�m�L0H�D����K����p��O��+!�Ŀ��XVC[{W��:�n&BS��EM�qrhr
�1B�A|<��b�->Us�����ɠb���}��HQ/� TV�*?\�����_x�'rP8Q��$g�vq[|�����T\m�n_��v"��s��t��/e��u-�f6I�s3F2�p� {�6}oi�O����b>t$���bh�8�^��L$k����rh'm�\Ӫ9~z���͡���-���c�ݍ�7�����2
�o��XS��v�:�- �l�cc(��IΥ�0��/�"��5�Ӭ�%B-O4{�+�)#rm��vHe1%[vm����p3��m�Q���ҼIJ]����@�C{�� �Ty297�PP7���h!���O�43�B��ŵ�����ʆ��I@ԁ/[�� UjC5/���g@���\S�<��=�d�R4\�H��Tr�(������w��C2�6����� ��U�2�����osw��9�0DLN���ؕS����EpgQΚ0�X���ʃs��G��ǯe��LG��t�N娳��Y4D�T0L��e���d�w�k��TL}:0����Ms�"�v�,���}�|���G�]���=�9�|f���71�>.��#�Y�fhƬ�y1& Mu�@����6oJ�|����bT�@��Z�sk`[֐����^0 Fÿ(� ��uW.��J
!ǧ��]�@=����yNP���Y��_y5@��:c��A`w�4({����U{�/��.�U�A�?�@Y�ޑɯX����X����T쟸�{���}�c���û�H�W�к��V�3/۰��`�p�e�	�,F��R�EՇ�Y�:���S&�� �	�P�k�_�e_���CO<�D��Xw[�'0蓽�}{W��	��@-��+N04�e�Y�sk��_R`'�O�"�P����W��&I	M`#1	���`ҥ�������+����`1�`�<;b��y�]�	P�8KB{7��'��y���:ƣ��w�4��N����'㣭{�o:m�� 򇧩�L���u�b�ߢ�U y�f�m���<# ��lQ�D�X��սG0]
���\,}s��%z3?�֥�2YrV�pTb����`?�U�p*�j���?���r���Q˽նu_���;�Y�D�����Q.��5���Iԏn�F�d{LZ
B�h7��D5Ce8���!n��b��)�T�=P����|������%h����N��x��`7���^��3򬤛�-Q�p��b�Z����j⫝̸��3B�iQ�@�3nH���o����
���&�t!��pF���=��5RZeys�U���+����}�[�^�B��d�����t ��l�^eVN����@�r\<�!� %C����o�	po}+��7�C�ձcD��Z�%���^�;����o���6��VF�Z���{i&��)G���yR� ��{��f�ν��ʨ?7�x�W������O�{�����	y�$�bj7��<��[��r��6i_�U$~&4�T���`�kPp���������l�l����FNCh��#+৴�s���-� �;��{�����F��N����y?�Wl"1�M���|����1Q"���5%�8�)��0��ӫ@���PX�h[H��� L�G�'2ݧC��ɻV�^����%|�Z/u��]�3�v�Rc���#��lʙ�?�g�`a�Y� ȘM;eؘDeIb��;P�-����%��&��w���Cf?ۤ�|���kb�����~VQ(��{�`�v��h�������K��Е�;�'�%�T�>`��0��a#�H���~-�/������Q
��"�P^k}����k�m|�x�s�\}-_`f9�l*,և�T�NW�R���%uM��Y%;p} �o!_QEәH)���E��,�k9� �ɪ����'���
%��k��"3�j�S�[h������f@�
�